// Amazon FPGA Hardware Development Kit
//
// Copyright Amazon.com, Inc. or its affiliates. All Rights Reserved.
// SPDX-License-Identifier: Apache-2.0
// Restricted NDA Material
// =============================================================================
`ifdef ECC_DIRECT_EN
 `ifndef ECC_ADDR_HI
  `define ECC_ADDR_HI 5000
 `endif
 `ifndef ECC_ADDR_LO
  `define ECC_ADDR_LO 4000
 `endif
`endif

`ifdef RND_ECC_EN
 `ifndef RND_ECC_WEIGHT
   `define RND_ECC_WEIGHT 50
 `endif
`endif
 
module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,

                 //NOTE TO CL DEVELOPERS: 
                 // The below two parameters should not be changed.
                 // Changing these parameters will cause place errors for DDR_A and DDR_D pins.
                 // When set to 1, they will ensure that DDR_A/D IO buffers are correctly instanced
                 parameter DDR_A_IO = 1, 
                 parameter DDR_D_IO = 1

)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   input[1:0] cl_sh_ddr_awburst[2:0],        //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[1:0] cl_sh_ddr_arburst[2:0],     //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lEbK/U+kt1+rj9V7CppSF38M4S99bZib0UAY2XaiLiYPFNJ1ap5uLGMOgZL4A1r6r5L60HNC7deu
lEQpMbiaOJ+9/XHEdM0oKmucKUL/49gjoAcezH6qEMKymTOrJAASf1/UhkQX5gpvaZq27AH7+mYC
Phj7XdkAnvZfGvPJMK3gsqdSg69iM69LHklQJ0+p5Uon6hqiSYzdUlTYrjwXfBzrymP9iWbSf6W3
VRRVUa/w8HkU3uN5k+fJi60b/NJFfxHA81yJYd0bhjHAWk+70RlA1RYUiqwdfpY+rlRleQU1/uJ7
qTvAz4wvSTC3xnP78ODFt0eq9Y5JkHeXAOqnmg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DJS1709GO5a1CijOn+o1lYceDh6tGAPqjd8QeO/8qiKZQkm5PvXeNr9FEgn5vRR22s2Ut4A8GbqJ
qQO8G3RxV9le4nVvya1DL+pjmHPCDskmZ7pMzOxfI9kF4vrU9RxRaRIZz90CtusVIH1SDYEdvRAC
rPtq2zex7IgP38+BeaE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Y+iVF4gwYrmMyAm428ks6WyeEmHDBdyH14ItNYcWPL+75ZpwLRXnlYFeZ621Y4rariKr0lTVQdUv
2CKGCWM7Ccw52eBPvaq1jvFMea5aJduRAgxy+z7VORC1Sv4d2O1mn7P9tP8mC4f0/URJpDIBRp91
4fYOJO5VWdtG28OoGoo=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
NbGzIU4MhhZccQa4o6dd/AgyjMS3djl4JW0Bw63MwoYVZn4930Agr4eJyTZaE15NBv3U5+PeKqPj
jexwt66LCA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 76112)
`pragma protect data_block
Pa+/Zrmm8H5eB4zwPXHCOimCvEqZerw9uO3RS3UB9ohSAX/6hEKG5qv2rxZJWebXPXJXi9MwX5ff
u1LWpCX+2/OWtnCRHlvYlYURTPtyiTOot7Arvn0/eaXXXovVHMPPw63U1Vyr42XSYK7v92xpzdbT
4SeAFMQyG0xWnhiwXJpV2DNFaxjy3JBlPB2etrUlUPoQUFeuZ0Ioxj4RiH+QHKwpGv5AuHsGdcNG
VA/sT1KzyFI9WDtNIGF1DF1vi1z6XwacwVzI0+qIgI13w1ck5CCu3IGR8LomEW93wngtlKPR81o9
p8SqwSVAGTbEOZ66RFThYjyPyqwvKxetVLashJVmZzoIMj4BkrRrx6pfdTj/TItCaxXvs9FPUGJl
lCzihxjyaL8waiwuKT9Ztu65NHqOCwadLJ1M+nLVZZwIvA5HSTSkUZNMsihWlCpMXrWwx4DPPZ7n
qKUVwLGyOmlzh/7MbJ+fNCIyeir1rgfn20U7RcoEq5B3kSKoDUbk47Ocs+om0d1Cf5E3Yjn+m+GY
iz6tgUrH2vSRpgDVoppurZR4gSBtwF9wTiBLw8vHpWg3/DoK3EC12EKJ+qK/9GquUbggDJycrfir
jqc5Vjpqya3uYpwUXA26D0jP2C4g/5X/R7x3ZK64i/8UzW1otm3/owO2k5ib3hU/BlBuCcNx+8gg
UBHbK+p+KVWXDSOrXW9xjfCWX/KeN9oFU3AGGLwS727yGDJ8Zvs9HBAPtgP2cugK4ys7a2XSEOca
l8CvTY7Ce8gI1Kxai3SegzZpz8w/BjOm/plH4jmMvBMXuGaU7M3lNN8ie4U/pkU9G8i3WR7pQPT/
Myz23z3HglucofmUYE3pDv+PtmFx11hDYAdpZfXu5JZPkbeyAOgzMWOUUbVyNKA3qBTVxK5frXWl
7r62c+mq76omaaxC2WBkRAMhvk9FihXCTQl7BVwf6/lA6PUDhg6PD9y5kdZjv+03CXA2NkXUoyey
0wSU2XSTaxiL+Rge2XlX0YmHf096SrhYBVnRNfy1/ZYIdvJ0jR8uXPsX5q5KeSc5kmcqHgsUQNN3
xMdUYsuY7ctlZ1Hos/FAI07Dkcf4k0+lR5iWfLCKhMBR8/rZ1DTK3K9yUX9//irTYwX0BzP/TjqQ
yWhyudeUCgBkRuQTxluRCIyxHLdN2PJrhVW0+abVyvKEtmDVq3AWHr2TXmK66BL5dD9tRbZCc0Yf
0msE852RwdC0AmXgwTv25SpJxJVhAzQx4IqdMJ1QdkQEd5k0eYiR1SbPkcuHlE7/bKZ3v2flRotk
wgzSZj9H5brUqHYgz/Y0qOIQuqKwlMQZRAhYd1L1XZJzbDR8eSupGU8qsbczulI7cUYe+Qm+QOVh
tD/2zVsewUeFMjvr2rLQONJoEiozhLe/O/tudTguADV49LF5S0+ICOx93K/CSMMyok7q3BvvtZ8C
ZeGsvWSFUU5wwPl80g14u3VCz+l2GuduqAXx1/zeONndTchFomFgWdo2FMkKcq6ajIJzTo3M1j8K
VVmgakLmvj6z5CJ8lAtei2tA+syuJWenb8pjiDwCSKBO/7GVWJxcGIoKYpkfj4CoynqsbLbP5VIP
MpCOYj9Phh5DW2wF1Ql78stw1JRi+heWuzmpzy63UEAInHYckiMh+m/6fH0WrHpBBNBUwzXvsD6e
9HkN8RwU3sUDYOn7WMnuZLVSo3xwiDCnexVPue511cBVaadz5vG9Q0ydxx9+Vt78JLnaeow3rSDs
sozsit3r2UemzpdxJ3V4Ut3Q4RAU5Ppqt3BNCQe0xz/nRrbqrex/DmYwewOHyo6jR5U81d3400zQ
YM4we5i+r0VIbjsMNIljNluVrlaf5JBwMrxbY0f1ko9T4v5f6ZemDagOMj08ljKcQFp4TO8H7I+B
bIUUfj7welIMf0yoHouhJ/9ONI5tGQmxSdn4Hq2YBS9yvHnEC5ZG5hkoV12Db74ZAHw3WSie1/Zv
wB+IQFtXtd5g26LZ9ssYweTr99eAIN0LBD+MB6uREtldb2FAeXw9uTEptdbG4S1JwUUOdPoX5JlQ
YebPTUsx+PyR3JOqaHKvmh8GEGl25dveiolQotPRkIOXNjN+6y7CT6U0VLAVwR4hEwFn2XzvfoIP
fYyTHIgXZeYGnwlTUvyqcLonAW1WP8wTMqWEnr+Xtopt3jLCsPIU5mfvXgwog4Z6t4Rr2g2yR0A9
REGAR76D8OnqKEyCZG2QX5y0SLC3atqMicOM6D0DVgEemtnCRC1XxzqP0t3uCZGtXlkMXlr/qf9F
ZdCYo/Pu0Ln+5+cmLNy4UMHM+LrJjT6jfVkIM8sJFOf4aw/BPJmlw1Mxjhmqy0DfHdoc+9tNUJsQ
OEPtzKdTqw7SX6v4w94Bq1gR4EAC0Z0EfyqOdzIlUhtEqFSsTKCDzeOHu/Q3HnXtF9GMGPvSnagm
b39XRVejkedJ5nqhzNEbk3wLtnANCsnoemueyc+5a6Seboo8srMhe+hl31ErqxTHtEyzdDtTRV97
sPr55WmvR5Qw2YSNdGdXbDfMxpdxM0U4L9wGN9M5lKEu0EK7aY1m73HVpU/VLz2oBbfzTeI6Mi33
X+kJ+27BIJPPa5a6Rdi+fITaSU6Lq43fT6UySW6OfBjw9kq3xax7jZmensXCOKl0PjxDPUtxPirc
gczc9VdVcyTUDnMqvpITq1G2ETkXCdlfL3R5pF5uaGIM4FCxFqd+7gvg1V4yPFHI4y20LiknLWCH
sHIPSqvdyGYwh8koXOnnBvD/myTwurtjzpaN29vuWrUqnMEEJS5efE43uZ4L7weHazufQ2uFt8sv
wKs/hGWdtPFqRRb8Z+YHnUePWMM76jbRoyQEaImgWURUiGYp4q2nrYTD6YHG5+uyJvbICca9sv1z
u6GWwrLt1VZHUNLoPuzusT99DAk3nQk7EPXrCAvV4nd0paYzHcJfk0o/Hr1FA60upOjOr+ZHvKiU
ccPq7iyKRLx5vnuKBgVoNNq9CxnBbL35Wnqsz0yo/UrzS3o+rz+b+8A3A8wV+pFpyFk6ih+drKG3
jZlU2VVpfB0tnoGyOJ+ZE1Lna2nnKz5gccBMbcAD08tG/vDu5KX1rW+8zpFDlg6qzgWg9k9aBn+1
ZPTY+8r4xR6nKNMVeH8vkVl2EcAhDTVkKP+k4raNRadRcoIF51vPwisgvgrdZZKI3Q5Mq8dFUsh5
RXq/NJTH4Fceh/C8+mdLvUhnbc8g2tXrPOh9Pe0enhO7tT3Ig83EJrrpUf46tWxO66lN/Y+QwjKf
WsBVtBZGwoubZzVHbX4NYe4gX6mdHAU7FU3Ul/YgR4I6B5ywqQOq8NMNUmWVQlvcZqHOi7cR8/Co
ph3eVsba0VxMfuFPQgZsdGeBA04jWiFJKpuRwUlW1bM0mlGuDZaj4D9CPh4cw7XEQbT6ccSVASzU
mH4gvmIReJJMjUbTFu9wh1vN3oPk07lmNL8UxR9m5BzRagDq6bURBqnXf/CT0ACdSf9AEEfqV1lv
8V88iWrvKOkHHspa5hUtKATJc1KhezdZdga3+mE9MaAjNp5E5sY4yC1oeCfoqK3OT5AwPg3lesva
E6pux0UUI2lw71kMuGsuhI2EjUVfIO2OSS0S/zV1Q90lCTpVMDDkdZJjCJrEHGQnuhRFOz94/4TF
IS/lpJDqrx+hoNxeJcd5o87zws3L0rw/io6nsQHoO70/+stgRGpzGFFHsNtmSGhPKw64WuQMdgnw
GNhByZ+9+Q3FzoOlJB79LuI+5a7kU1IKCWIULEGNnw/FXAl26Ki448lnv/CQthBMvIV8YyvvoMXn
rO0t6jKZObLErLiWmh/G4je3TSJPa8T6ruVjWghAa2u4iCqKVmbvIQ/7pSxTCVdqZQBaxuKsRiQ9
iia/qNDsGAbZDk8c5v6fyx9YiLweNjKV3UdSdGb39cnyFKrzRwjPelHCaa2Ti/hEM8Lq5dtlsENC
dyy6ti9sWrRWD3dTiCaV0gV+2fUUW2vQoFiCo6zMA+pQDAHBvaLpnXVEcePJMIJyhg23tXpwrXZm
VvId4Eic72QJNW3tTzSJIeIEiIXkyCol1HQ/KH+wBFCkQFMVvnSU4Vgq770a3yosTie69N84eBJd
MjxpgtRqaLvON9jeRPLWQwuwVd5PEpUPu8BHG7gfPN1AlATL1Lvrg/uicnikTtNui9puPCJ0HPw1
HKI+QsuNsQj9fDyvtdTe5dp+a87IYYWQBIjxs5hywW47MZlp6ogjwL0hSFsJS98NFGjMO6Fm6ZZc
5u8z1UOIrzi208KSdBMMyhau6qZ7eTYVjqD/1y60UjAg4xfGXk95nPsMEBDR2GWzJ0ygEihjpHOg
st33lXxsV4wY/lN4LQ4C79Ll7AV76WAv2vZ4VBon/dbd8+Yl40S4vLvqEC69WtSMkeAqPyEndltp
MqQqI5u/TT3RrXfiusRC5dzPhCwPqsnCc7A+1pK6lY562827sBmlstTzTdjIWwT2JpQ1tBl1z1A/
vYi8Gfo9O3VYk/yCdglceNQr9isRLDceGU7cZ195typCs2zpnWvfgEQCikVdChTeIHoU5GUyv93M
kYfFU14k3ErWEyi7lh7vUES2AaSqZ585EM2BxpTONvDGi8Od3HARRa+Kvi2QktLSFf8IPDXK/TKi
fkq/lW9vG1jciZz7MJPVDQDPnP6BHERcirtWDTlWaiACOFZbvsrO0NiPRhpnTa56NhSNY1eObB+U
BighnFTqGAAewj86JjkUjLrf8vekKBQcjvvZHiS0lt7AsWmt6YslrK/uVGKKVIdThZDnEyB3DGBO
/VWiR/4IA+Ayr4vv1dNb9ycQgAqRCQT4fcZf8MCynggA6S4iQ9hhAT/bh8x3xUGQMI5hZ/DpIVzn
+KYlS1pVXowewa5KjXbymXvYJL+5ruQFtKiH4wMjFrD2t1syizEwkpnQTD03meAnq/53tcdST7MT
MtQ2NVJyb4PcqebDKiNI3i19bvoU+RfsJt38XQJlrz3BE8lv4Vqon7BiSE5a3coWsjNUOZjUNMDx
N4o5m8/qcclS+2NqmeXa3fdYAt3kV9v2Sx7ucL8PLD+y/WQqgESTzDXMBIzfiq7bb9a9WkCOp7cj
HC1R7DZzJsw4SzxBEmdyy8tw2Mnj+2iK19WZ3EnxGhX7RY272IsHOlQsMzlSlTKBZADwDiEU2sZ+
mMSrT6XhcnxnGYDQSYKj5hKTMwgx3NMXQPDGKAofsJfobU2/ptHr7sc2FlBq942HFyT9Xhlt3xUR
EvzbbAItWCQNic1aLEQulGbY/FafXQRppaToxAz8AT360l8+nsfTKatvEwEkFHVC91rGlwxsx26p
PVf5rpS/NFWdtgYPfw2Mg6lPSbNvlDtbopMJnNEsyuGYMDfaHQzZFOFJikcLXTQVYIzESqG4eu3n
SwSC/E3xwnsx76HZZoONOPV/wRdkcO1t5FQiFpeWLrNft0SQSthmwUbsEF9gUY7qRPIVH8jJqOAN
dujtbrvXqWr11dUf6oDv8Y3amTis4vpKHyKOD/SpYYxzUSF3UgWbz4HGaCm+Y7dRjxMmvI54ruLz
1wvpMPWVOHBhXIAORt4+7oznrW8JuBhQ03AoaE43NY4+spayy+rysX+n+gc0CegxAnGi50lrm/Cl
KYD/pFK4cOd2w7+2apiQDBSwvQrMpDcCjgonpHYy01roXt12RZKsyq7XjJgKtPrW+2UBSzTJagtu
etXbomyiQiCC6MWyaxc3X/AlHKatfh2DiMQZ/kiKRvBAAA4X2tSaF9xGFK0pVklWrZbSrkA91HEW
dFN2RBahY340pDNMy/evmLOZQiKwgVchX81zVcCcsnUrcekEMXzroniOllG7Uyu7UGQzclfYBn7d
pSeU4aZfXg6m/szWwqgSkpUEo9MXxxVM9+EOfSrJJbrTHi06xRd900mtL658MJeAdwVhsnqilCmL
HC0OE3QDr9ISgme+bFyUXWkY7XJVlQ3gyFpXYmWbqcPek6yhK7Xo00U9sGIDFMI9CwNQb5eKI24A
CuDdS4aMwk3b7UaGO7XatP0vf/pAHD43udE8x4xPAdqH5CNtJsbj5qeNbAlvY0G7h1Pm+arHlrFl
d2h507Qkcj3zZcAdjf0gFYRDP6Ihbznh6WCk2V8TWcRHw09LqtIqrtlGZIjXPk0ujmcgOi2D7upo
6Q69VR6RucP/V5gPa7WbFIkyIuffFW9EWIYvTYT7Uyk9Mzhu+3Hij/UOJrlPy5Mv72xFdEhSVySM
Uj26VdTLfLaMI2uel1prBjzPup7o/0FRre6Dj3M7GTJwKZfZie9jb8XAiYJTZL2fM/phA2dWCX2a
e5DgiYwruFInirQ7l2Mjcdvq4suwNeGUlOWSbX5S+7lZ28GiHwDSvylp0Cxu1F9MXx0kFOuZIawO
7ccq+illmj4GCIUnfKWzkxyr7NoyTE2s2RdFyO+UkDj7zb0/3Lxmd/TUNqLGQ5TCLjsa7Ik13AcO
4dnoM5XeAGAdVlmMdOMMeSnrefUzeoTagcWnkfiCmEDk9P6INYeslJiXGM+ruTsRoAcODxyZ8e6E
vzcaLQ1tm1Jq4MWbn7iml50Z1aPvdjtBvVjgvNr7iQ2pAEEixsSgA2Jnx8NwSKlArs11C2c1PFA3
La+/wb3fuHNSeO1GxxgyvYiSegbafqHf7J+GWt6xhH9/rBSFZ5EXji/v+f2KvjS1EmmR9cNAjKEf
6J3q10DusblWq/RwgOJcMxIWxi5+pH4YJLusE5++H3F9mHaxk/FRHu+76WJcM0UtIjhBwcj+EBVy
joGrq2n6WvX/dbpzU4oamE2cX5H8hlGDQRF8zXQabvTGpvLmJYR2RPueRbmHmwtYXHlIMFF+sGKX
iar8hf3IFGKIWStuvRM19Ay+T7pG8pgtDyGbeFyuMd20a+RamlfCwXFXRjSqDuI8R+niqSJSe16m
bmIdAURT+8BmcJBB9/UxwmsDu/U32mZOUK+WFMQUUzL3XPQqjSWmTMSR8TYHb3BwGXeau38yBDYC
kTQ3PxLpcJJB0xxtUYtgQ0SCYAtXoTz3dtpXMf7ybCqhQ1NYri+sf5zC+XDcjohCJEKR4GuLBOiX
1BYOoQQqthu3ZdIP3+DAoXiWUSULPplkToIbhJrF0BL3ief6qFZgNx0BX8Sn6GIeRpW6FCoKeGt4
EhXK/kpTizavKdJuwidsXDf8BqQFlXU/bCdX/7UBTBvBmnWzdSUoeofYcJ2h7g3UjcO/DDQK1bd7
HE5sOrQ6YWkEHakYEFQvxAIJuJOFBqF2hylwNZiynf55bT0YxVgRVdk+K4O0ERPb9oqVorPDtsxx
SKKG/APYBeydaCMO891J26MiA9lWUyk8dukQyDlphhojnO/GfBrGRkL9cF1FCXHDp8Gxjknkduft
96ygiblMxPjIsaPKMD25OChSgOqQIRsAepxIkNeOg3l9RVdkZM2Kn8B2fkWcYkYnGiePSHBOOEWL
4rd/4rqizg2NDf1D3SVXzD9NtGfFtyCM/wtL1CfvV6IrX6KGH2z2j4b+ubdHSj/M4P34XDrFiYY9
HoUuGMPG8mVZwiQCIJdQJAyiEJhaop24nwqTAU362knn76QZ69H/j+J91fnaRl7P36MAYp0TdwLk
/M0VYqLbdu3psktwFcToZVX68sjT6Ir1lKPKBw9auAF/ZILbnZx8elLFKltt3Wb8PDyxLoCpRxGK
X0u7YUO3qUcMgceICeJ9/rCbyhF69cUuv76cNUpVKG6W4gMBiaSyvnZCCHwiYJXRr2Axqb7KHO44
AfhdihcL2EiyRkS6aqxYPtcUw+dk7gsALMrDROhMk/d/yqDzvijknkc8jxLF+f1Dyo5mqmH4V2O3
MQ9ZDg2m74Mr39iiWQWNpXkkyUfSnDXWLS0F/lEDuJi499Bo4RlkvSd/a+ehMaZ9mL29qtqK7Y5K
K+AVoI5XUL6SEPNHd2fIQa34IRgFYQSW+qRsuKhhw+rdi9W6BytXajJBeYMdS209xCCXQ6SnAyIm
1NHq0U/Rxdfrve9d7CKqYz5GZmRiW8IRE9KZg0XMT+IhpOnZLnOMwg3QJC8z5nUr5PbJqt4FztM0
n6RsbWlobA/p7eyCzX0hCEN9WV9xYrXARtlLYXhjhM2GcU5K81UCDmirNgSG8pQJusJ75dS9J9eA
j0lZSm3Rrz8qF5jCf0I9HPLDr0pYq2vSjO/42Lucv/ZWAfYc1fjr3sman6Rt8rRTx6+oREqsv8iM
oAQ22UL+AzothLNzohQdVgiHEnlRjetszlsltVhzEvQAGFnw/SM0x66/54Kgw/sYbNgzswkc/uhR
0Fl6O//Xn7FKkJKGLVsfEUVHlT85u6XIKNE1Tt/dipdYqD4Q3RBFuFmbPvm+Q163P7muVP+NYwvY
9A2Vzz6ZS442vbAY9DvJ/3OxOJY+P/mWLYmXKJ3GBP2snGgHpU0LlOB2H+fgGdy0+RCYCyrkglQB
JAoIYU+tLvEji4UeCwnGElBfMPU2s6XjMAKXz9h9heeF2y1FJor5LMspf5sohYsKvi7i/i3bUl9f
1YeedW+olRShUcKLPmFgtt//bxZ+2l0JUARECsn5HGQwri7EcwRHPFcklOHHf6Fk3KB8S7OtMkJ8
jZ//Z0TPstbeokUUphd49xGoLEM0c6LivOdIf5b+6eSJo/ZLVf4T01bIRdWWDErnYDt+D81C/5TX
H6bea8G8EOkD18TOL8GXOcE8rD5pPJXt3vr6HtoytfwSm/2aOjiipa1DEHfC2TTjRODK6lqZJ18V
6wo7/+wR6JFhgTU3mrHuP+gPHzIOB/7CMjECsCJqLR0BzcIfQQe1ESTzVrDOx1udDm8YZlXIspyU
ns02bROtasKapvKhPdT53jXRWltd7f1udhxsn2ZBh6ePkw2iza6RGSqcYdPmzbBgDw8Mevav8cVU
htGROTz/9NRXCXFgq6xayDQSmz4t2pvlYiTXE0wPQVMELXQbYbEqAVPexubHr8wWlPooyG8WCctT
R1MKZXl0gfM8z0wDOwIv1G1kCewTz0IDucawgBkfG7eMfyxquldK+03xP+HWxFQTdBqVEmlBwap7
FtIKJiycrkC/xBbfuUo3qVGUWLsti2A0utu9zOrD+ULlIHSyq0nyaDLwzDunHp4IMnR4YWWp3l2L
0k2qYDhG6Xdv8bLmLQw+1hwiNC3q2fVAIMaLcrRYiSmrVlK9LkwGuuoqLJ5FQXZTadXiedRnxpmg
U4qrbmoJB+IvWZjIGuw1espcSPA5KurGwhPgje7amFaDJCyO4HgodBk1TxIIv+h7fK2qCAMEubXo
+mKXpiwsZRyy4kVT7auIKkPB3Q3JSC0qeMxRJ5w63xG/QqV/681VFBycan/WnUv6q5wiIG9QqVON
1KXkg4YmyGKAQuDr6rPSEUqOSFtmZKuLbNs4T84WLfpSFCJTn+pHl1/+vf1Gxysd0THLRXgK8r5o
sNk3RuHWOQ+1DxOCk8qPuEif3HLzofqV4rMu+M6Srl4VQWE3OuFPk1uJappLUBghXcMf1Jfd5rGG
3fDCDPOMoBQOK7Tus0r2EKP2d4s8KWY3zMzKw7xIxgCu7GUeNQMzmPK/Umgg77MOxEdLUp4FnWwV
fg6Hi0Usl4l0rUCZWTSub5ySCmHD3GdkJSmGrp/zJ80d0OPn+5mzD5W4+YvjOoZAGfLfex6H1WW5
3DjqwgqlIfk22X/T1FAX/Mu7ypGuEW2OdY9QutDHKof+Dg+JyJSCtOv/zA2AMTEYHR2kjqGmy+c3
FiN8SG+Oh/QwNDmkwoC04IukXnxU7mBxN0poZLGfYrmaOWVsowEkEVuABXmkalQL5OHiWj346Hk2
hYyLCUddaOlQYkW2RBiWwTEweZaZi53BTT6TGjggLq83fhkmRVrqInnIl0h29ne5wHqn9hxdBrXR
b+JLYnNDlDA6HjA3RUd5cNFGfVzBadR2QTo63ozFuX0W67H1/UizIs4ZliNBysIaSSxNKpunp5La
0wCHzqEkHZ96gUz1CdOo1tXyvy5m0eQpl8LPk47yj/n23fx+DJ27BCRgKerQTOQ+6O1LjCHGR8y2
HvUbYd/pyNBC6N1JE90jG3PW7Sz/4cHLVPUEjhVFxgwYDUl+zcf0GJ/oh7QZSHalSZ3LuVSRlQ0S
+tfs3dKILUYPnrntptdaz9uW2mLu68lWxWgAxD/IFp89JuNaUQXw+Crw5fcFPCp1V34CzgATgygB
urnF39cLC7PRT6uS4hhXuJqBQ2Salg497gqL33OmYuECU2k4dKcOWMpCOLI7TDJENdL6GdN4Gh+x
nNpOG07tUPfEfNI7cZs9hzGl2c/HU4XJqLZ02DrS2Bn1mbOMbcpoDBkPnHF+ANqpLB3xPJTCMvDc
l4XwZYNPC9YqBVomyMH0GOMAo7XcBJGAQrBGpI6BEe34q4egSk2PB03pAGvXgFGmmqmADuFAxIu0
NxMRvz/bjEk+5LxHKMM+T+HoU6k6TRlEdkznYVZnUefOg/5FEXBchohGazWnXOrRa3PqBI4Ygzd3
qOJM/SyPxWzBb8kR4QdJ+nOcgV+uLTF0PkOjyVO8Hg6e+2+Q7X7Cj4x71GMfxckkXNmUUJ83j6E/
MWD/boHENozRkTlTn33bOztmF7TyA6KMW4FSNOHyNi+E+Jq9gPHWz0pEkGGm8hdlbSIMxdIHu/KP
zIx6bnjDQvOtkvmQqkyX8Sa9NRiQIqsviFGCcW1eJVA4ZrTHzp2KXUMBOgbBsXm4yhlvg3iTUyht
EBn/IcHgBzPQGoYS+9aEIhiV9szMyENzqpNzIj0Og1Om1KG6gWqaQ22bvB2yVqLhDu83uCcTpdMS
/wEUqcvdbxV6RGa+zZg8D9p7v2mzuGBjowJ0jQyZdTtINQ2Wp+xDbm+HT8SkYmGMLjmbgdtXNtFV
HsHnILWY+EaKJJ5cpUhmPUFEYp4WowT/H3rG597H6pxIx9fm4Bu6SNRkbm0yc1LIvqBrUkSD0gOt
2atqFvAkUB+jNPJu86LxI39NaOUmILCwn/q04vD967TnXRjJUQABcyckIvsJIIoNXyCEa3lrlZRR
9Z/qhRYF3wK9xFjOxnj5uYir7ug4iw/UGoknCmYC64x0h3xyJigQKS7NN85j/S90R0PM3NXVqsws
yQNUU6AT12VFIBOoBElR5KvOQp8zI/56hrmBkch3kJBdGLbFIEYVH8+CKGtLTb9XwkGv3GCEH5WV
wcYFm2A+hZoUHSibxW0Qf8L7QAsxZDKMaXXc8EmNw7z3s7LEZdhmyaHD/CzxmCQjBgbMLie/YqAE
wvyRl73lpDSiWakKcxeF75z5wG+He6E8YKa0xxIG3dAJBE1aSNcPIZyQWYx0GQ0ioOY5Rixwu2wH
g4RXmvUo2v2ukka/MNJDMQThblu6Vtk4bO5zeuYFr8nWHNuyjrFgxsNL9JmMjEQOh2woXRQDcfHK
zDBvREaE60QtI05R3Vvmi2Yo7EjUWL/NWwjG4hOU48x3JVWWVwlFrUapKMprS21QZ01zaWb9GM87
LaZWyigjbfUTsyWj2nTEfPXOdkMz0J5Wl2cVne7TN8jlcEdJ99PqDWvLMXQMia0Gcaoi7u0UWetj
AQ/S5IHNSfgXngeMN4EzDk5eykkXOe0NCBvkQo/6q69G7BbJZNkTt4d+TUzYGGGnYUhQW28Pnxwv
xs4gfji3out7holY9+VZ7YmAGXRSsC4h0kbN7ns+FgFtJelNf5N4P3Mi0vR7SL9tdRC8YmJR1pTE
DUNoi38xTQvNR0aywFmP4rsvxOVwHVz4a4qOgXUnQ2RTJGrSsCTf8uB7zKLMhz234/L8FYYURue3
JxqSj8bYbYv//kdbHsniKHyUOFWIoJqYnVBDTfYXKp88dhCjTOjBrcAYCIoDW1R5AqIOXVrzhKaX
qQZ8HPehNmW9gdxI+5L93lav14SrOG7NOHOnqsLEoHDvlkBlXHLs54p/YW7fSuY65UelVPiQjdDm
d9xESz94YuO52YsDpCFc92P8dWravpzwNE5fuMiD9uqOeBK5WuCAgqzPJeaRkulhX49y4Z7TG7Ik
WvInIZfiNWn+Chi1K21qq3LDh1kByfB9nIquwhJnYhrPaFBZ8z2fGAh4cp6MEID672+2KxFqGi+Q
qCZquJc2GfWVxSyiIY1uzCafQVm8OjtZJDvwyX2j8u2zQoXcUjHn+pL1WaOHbK0PfKauMsuQ85UT
NLmSyFwfLRflpQjJvnFzjKLGdaxVV9lkupzh7XMnhlrVa9U7BjWJ18mfGMzyWAzhqhl4Qi5ZMwLQ
e3zdFBYDSqhbCIQwXxKCQ7LRuvOVr0XlXrbtMFStlvdXDhe8VID5/1O0N0Gdb7jTkjp719NiBdgA
eFE9EHYe7KGQ0KE43XMJ6PPS+0TnVOK9gJ5ekgggZ8t9uWsnX1yJXwiae2O+QsCbwW4e0N/UDzVC
6BRzi4YPS8HDC0jduJrNSmSBzGpeHgmuNSQFuohWfevlNX5hnAtyT2MbZ9SGif8VmzcBtHZLbJo6
QlGoJOha+n3TUYCccMNwh5VxMLprYxrWojN1qhL/buQGd3f5SZ6qRTLiYIAnx1/0rssEfwVDU2Kt
JST0eSGAPkfj1RgBslzgbmyNacskdP9UAQpfmeRl6Y4lS7AmP4C+E4xi4VZOcJ4D2aJ7uHnvZEce
rb9WgMvvs7JXOZ/IRs54EIhS/VATiGr7gK71H33+nO6+ARD1+e0t6Jquse2wR31VGTrm8xjDuYZG
6mFy0Dt6qqEcG3ND62J89VQayP4cEM3Axe440E7iuFALfMt0uT9QSaTEAiEHB75DgXK2Ykeh1lIz
tuFutOvbCu/5/rFXc7Mlfk40Uw3FHCDtm3oCivDg3v1KeEg643TmJ5dCRPCw0bycJ9NjkKvAE9Te
lbEIaBUxjRWhKmaWWI8X7Uh0k7L2l3o56kaQm5Y8Voi0OMql1+R1D/x1sfrtPmMW7/WJ6vjODlRa
HfTbXneC/nv1JumfacboWhMIAso+qT3kpfH0fngysHN5CC8k/FXaZrsGJ8A8XsQQQNgydBVBJA6I
3g2xiqy+vh2ybGu/59rkhX78Rn5wYRvjZok/fPdluQJb/9kkYUX2Ay5gaTxXm37VgK71d+VnEDMt
L/luciN/x2xlhMZAxEVZI1XW725uMkoW+tMu6x18yD573a4H21otiMWZK7n1m4XbxIakiQ7QAYsg
tCZZT6UkJZztUcF7PY5eNnytqctAow80nqD1PmyZXBo+36v4fNn7zyP6wdlyXuDCp50OLeE6hF40
YRxpLMyUbpLw8LRN5FXwDp9ELXWVlvklhV2yveUYmkWv/XKki+PvDZaUS/w+pKIn5md7fKbBkUOj
NJRDDM0PYjOpZ0xNYlpGOwNEK2w+qxOC3z6zV9uX/TYsIntnC7/NrSJtUFcpM9845OXIgMJEbYCH
5NH0a+liBZPWUjklXsqglhYEYdYekhnXV0hx/7pURr/LYOlBeLHijTxKnRqM3kAY70walnTv7EVO
uBccSbNWAhH43EbiHRu/GgGgs6jaZM7DZNXfxnUVESZybcNC+Y1OCwKIr80NIdHqNzsrpBxMlcAy
XU36KIQqRk+boM3DImhm9X/rHUu3YE9T1LerV1y9YgQCDf6wR4jUgiXra3z2L4Uirj+cOrbqRMBo
Vdg5bCFEnfT4nOQ0wR7aMsO7uGjNIebaNneVvt0/rx0VtwPo+9wxJBtL9iwEf2HSxGhaQR6lYYie
n24qbbPDhRNl+7luXjGVw8NJaiLs/kPNTX0OiOgj+TXbiwytCarD8gRHzZB8gG2RowRl7cqMYkQ1
JvRQ2xjKYV2OJjNnYbtsrrOFpkAYPdSLFZ5CQmWM1da0ruVoI37i2qviCEij/ymsxJ0hQKCm6SFk
clroHI6nGct8G5gY4h/NmC3zF7I0hOpSg41mNeFv5BqFNHXq2RYPuXT7k5s59d0ON3/OO5nR7qyR
6HTdr3mshp3XHujlDLnriWZgY0UhEe8arSP8qNj8bLRnJyxPj2aG24iM5ySn3uwM8MRXitAJL8BT
IUbZM1NWjvsjZO0DIQWwxvtCWn/C/CeKxdwLl2vzERJdBrDpir4GSUsoJXSaoicfVRXmANszcQQr
qDmBC02J9q0xuiDX6rrrccS5SzV0PiONjZTB2aSZYbjl1a86BnfgtsQ1LyWeUOZyiDJ27UMV+ffa
HQFdxj1Yhtqyq+Q/0nDWQLjiHRTstdDFI3qynE+8nDeOTxcvUc9FlyRPEo90D0V4fN/7PjWnd5T9
gATFWuCkTQThR97OLdNynKnoBsIAsriIN/7Lfqwqd2V64waQdPgQZyMvnMdlaV2EHS8LI8gF9Kcs
nzAscG4UPT3awwnixE9KMUBx7/vNpFneXxfQpaZaGQRQo6UQZ9jutL5lVe5sU19D6jpaWAz5vhnH
S6Yhus5ilJhd006cP+u8avA9YCDm+oe14nTpnmGX2w725zcWKbgzb1KyfLo5Ek5w7F1K86r0TEpY
0sm/rmwTOx8esIc9cCVvX5c9ZO8KvfkjT9MIhF5FKnTLjIos5sIkNEhQ0WfbsTTy9kIaFS3uby7S
jZoP+1sWuhYqPPwCxkYFr9LumPB9Z0sNJEktuBm0OmZndRuNoMs52VEl6sdCtjW+FAN98Eij4IIi
atUiuPb+15i0bPMx8hDvWiia4nBfP8gcSXXLI8qHoE9HKtc5U1rtKfBhDdSY6HWpzCRqLbv9/EYO
87+SKwGCCizhBp5cEbzSRPK3HhtrmiNTI1r1sAQGCDk1OOJxdiStlaWv56KBP2vnQ8KYkX61aWit
mu4xFD9G0UKqe/ttJbQQRfxpkGawmw2DBE9t+kDyoQtyz6Oms6BpEn1IfB17BEDLzzyV4pPOkDSm
zo4lAvtmRf/p+nSkMBHIpJZWSRzXQ3ikYiL64WRrnBb/32eOFrTUG+f0eT8axTlgM83AG2cwZ96H
rFEjvIa3sPJQRfhcWy4fKf9GiQjFUmcl/auYxNHrQUP92XkJyXR6u+zytniRn06CAYyTrX3z6MXY
vB5ONECkEJwnwUSRFSC95DEzTI3xQk9+7PvVP0iR+rLPITsC1jABJhe/XHVyMf5Ed+Et3MkS3fNw
fKizsxByy0t15Jtt1lJw6I2Wl4Y+b7vARf/piCIShy+Btkc45hEmsYed164NATaZl26+Y+dlE7QY
PW/IKA3nD5ukMisd/aqCaFmtUkax+gE9h/wYLbG56qnSdhb9MAvcG/6PxIMPa2oHlwZscil4kdLd
str+VfCyGywHP8OUhfEW/Ex1FS6xjvVaW+B1fvhOUDiTHdPgdocn2DVTAqhbt68LMbj3k2rYlhzu
Xgh/UO1vX4nyN/xaauB8P9hVVbiGTWXKxLQn0drwZjyL/Z0ubOY+ZwgaJw1z9MH+iw8adz6DvWEg
1kj8TratPZVrm5g3vkOWj7N1rTP+urimgWr5bpxCKRV6m5GbA2Lr4vzYWg6XZ+tJll3n8HJgc9TH
/Mh5oB7h6CIIuPioc5KxUx+r916L74XzqX5o/qLtThLOAZtiCBwQBWIKpVzormadTGC+1HHYwnc2
rncEwyABRM3dRv6BgaWIcpVPPgnpcz15l70rcifztMZYzXCNQgFzlOioOnEwHSfAr0mABGnCdydB
eu+xTamrV7mjlB+hlVksXowsmfKVzGUyy8Z8CodujJnSBay9dRIZVN5wuk950zucrKnpzGifKwmV
YmqtDdc0IS3FSYjwxDeH7E1FFV29OCexbmpNNmLdrtLrJXWTJgITF6yD64dWZE5RaYSdb8sQdAC+
SYjmKtjIMaynzS8SsfIlTAa5cw4C5xO8QozA5Wtjd9ZGCe8sJmTJ8kHUNcbC5k/wR9N/v7txHVQi
0hCC409vds6aVM4D0EpeZ4cWWzLiyb/fC9soLR1mwiAOOZpJ6/ZHW8xQUPM5jV4GCNFKGcETGpOb
wk/ORO9x5RbIo9KowCSvcUpy+xEC67WR2uBK/XQJNKR3zzvk64wYSsUNeSR20J5dxbe+BZteuTGJ
nz9VZrQqyQAGPECRZnoI/9JCygYuI3Vw55s0en/PogDAXj4JCc/Q1uL9f37yX3L5ymLAkxMINb93
zuVcBt9lFhgm3APZU9qGa4NtGSlyJ9fWRyvBaVK70i88ST7jE+k4DSYE4w1LRh5AP2erUWSxtqDN
23jWafrWK6nxkq0vMCJTA9VhRmXhPNh2rdn8OZOi6C7KF/V/ro0zXa959UVguzR+80UA3t7iy1HN
yFhUWEqRO2+Erx8jE8/vCbHTaupLhrXhUTkQm2rXmFfxNYV9BQcoL7AEj+/NZpFfxFh4+K8EF2n3
Mc8KncjwIid3Hb0UOX+vqiFgdW+agKO4Kz1VCbjrn6T5XA5cwWt2dNBJrLn0UpW3pmYqpJnl8PJq
nTcOgEK14J22ZRCQ4NUDMO0Qe8XiNJSWjFa/UBeRFVwLMwiE+DY3CfYZKALeoRRzOq9kX+ZRB7mp
ZJsZTXAogno88vGUqhFTjEtKnzNG+gQ9Ax6rfQtRvxuMlsRu+XuU4EBlxguWHwCO5UE51F+rjVtG
DBnkEFB5xFqIkoGcrB4rbDQ5khPUiaon3WPZAG0SAaV+svdkbYVpFbELb2Ysz3g4eIGjLFAd63B7
iWqs2xAAjQaNaLHGQassy3nN5zSgAwoxCSTkken2i4xS0VAQXvBSr1LB32jMmv9YXq3FgY9qOs5t
T/5LNamZEmN4yazNanq/sa6LyJ4V9w10qYxdym4CannzFmYoSbIR6okjazhd/YgbiO4uBF1aReW1
2aP/YNlh8TVLjCP23jWKNEzjwNoRAbVLqYR9yfskoFpO6JHV4xkxV8ZYlbvz2Y6MC5eZEYyiU1Qb
iM7XXEWS3hSGuy8NN4yznUbilbHDOLW6Hecdli0S/QJyq4EFEAjbZwgVKpDRzqoqVVwDJ4xdQT88
tgwrxFcMImNt2kdjFnoNLn3JrHIufvnMkMuk8FIXPGvCNCna5z9W/+8UI6HqIRrhz6+rSAyKGB4h
remoPjXUg3BVzMVxmtBSQ7k9KruLKcvg+5JpNQqU5xiAENHIfwqDUNaOLD2UkKPDceZjQMAW3iYf
RDAKgN2otFJgkRtY3jRnOKjwJKJXnfWvjeB8WW7DWC+mEGJcPZtnkuLCIOnOC+GYOoaVvktGqMbz
1Cc2lw6ABC9S5g1k/za0ebJW9VnqGp2DGcqogVMeFuuk7ECcfhzcKV6A4cuENMBT7d1LZiUAwEdC
BNWMHEknIy3+F00rv7A7hrP01e4jccaYt/kb/seRA5AWVqQCLU25W0NjmUYq/tLgYx8QnWNH8rZF
2tm5W7c7mXK8FOe0ZiADc1C+Z+AJDOpizghT6dS9d3vPfa5SF2r4pZwR6dFeiVFVDNkPIq1NfiU7
YPEtRdXCK9hW95Hu7u1igP9PQCmOMy3uSp410JeV7pSiVEPrCKixE0BAr9+cq03VL1yH3GmQsZXx
Zsqh8Hh8BCPEhBOgeWg7xM9Kcgm9Kfs1EV/vzJEfizyI95jtKSAAKoF6ogoHAaPiKC2lvYWpwRfe
LtT4zs7KtRdTb7jHkjrlonOvAI/2lIQY9Eh0QBGUEeKpocZn3tDBRehdSljJENPJh0pQzjtw+bEP
RUpOar431RxjwDBB31aRNKRqIqd1Pw5cxANKOihaF0WgfyP3pkqqXfRIup5x5xcQ23956pi8LLZl
BygFSgaWCVwmqwhxwLelOSlcIh3G5Ghz4c9hz+LYSPkgoBppS69VkHX/anjbvr5tYRIxGeNU0Nkn
Z2/W8x+OcWKp5FooFlwslZYbmcuhE+wxqJqi1JBzbCTLQodBgF323lRgfgun75h3VKc/QRPq7Rtd
ByxzYoaQKDw+eOZGfPc26N1hE+oNkyCUTc3BBy2eDYUkwE3kmCkQyrDsmi+gS6V6Rkm4faBLFbXd
fXtyFw0uhBc4tHJAb95ZfyMSNAx0EjQR2d0+1ZDjGizd3pKEfKDcAw+Bnjuad6UXgGMgRKR1071U
VJYMYZor8pSDP9yHSUAn9rIGKjsLEgZQnzE5VZ4wn12wUeXFVpcUmUdggFqfNQ5IHGnLWZtrLVPQ
IKnxy8anWR+qeh+D9kO3ulwY9MWXdOaF4v3F0GqvR4ia+1+cUOlqZ1OTAMra4AhsNibiElrg7qfb
wsySKfA5TZiiYfy6fdDRnVzFuhif2IXc6jBl5HjZnlG+S7icBo0y+qkZfPAWbPvbm5Kpiq4KzhHz
Zdz3Hjcqr9zfBsrzO+mC81apZvg4VAK4+ZcCPhzSaK19jF+oqEbNRAtUHRQ6BwVu4kNyh61ZPtdR
ee44J96Soi0SeDCA+xyfiAmaP2LLWYhcwwwMHKYqaDID/0s4azuBDdXp0eINmFAcCTPv0trARGJY
4N/1a68uV1LLzA6RlYf8aJjWYmO+5KxbaD4aL8gW7BtJq1SsECmvK+8autpOW8XdhK4Z8hI5qe6M
zEyKer6SkU3BjD/Gx+2om1hypJjdtCkfajqBF7NobCVDudq+broVsUqqjuR7jrq/mbDIQbQZqysB
1SA9ONP0h/ZGCwYwqijykNBiWd7aKyhCPH1ZUgiNLKJw4YYeV3kkuhUun/ltA1zHLK3aJo4tLSIy
fNquOlvnSseh9WMAmLMD4KzhTYnl23Br4ts/picJzak5ITmQvOR4XPKfzUaetAHGQ/7D+be5ePL7
UzmEfRTKTr/x5RR97ArpuwxjRNJNqkPB8PQ9wQDVHhmed7bM3TtPhzmyPpTVTujzW2QdXULccbf8
tcTwg/Q6Ep527GAOOx6AQ/vww0ZIvZhOJA1uJMkPIfnWMSAViS/VojA4BEHvuZohZaiAtAJ5fYkx
zpYi8vDCiQBox6+LY+YZfytTYt68TMHT7FphuHiPKVDlG7kQoQ/HFo1uamrEBR8oYqjvPloZ3R/A
SNFA+0liTMQiyEiHWiVOL8KGAqeBOA1Ov//J/JCjYlkCfmJbl2N4lWmd/y0RHFwRZivUONyLudeT
Az/x9hBzM+p+X96aCMbyYg6gqCJAAmR6k1fb0yCC6YxRwCjsgGAwsjynBQHhp0irIP11uh32n+QB
KK5rbOhtE/WbyGNH+63DJO8/SHLW2AkHRx5ZG+YIjA0+c3nKli33ilTb7BTuvLzVJRi5F1Vu48iM
W3ghW5HNC9igo40b24BLTp1JlOrOA7UNDXgwH1CnLN5ML6bTbM0VV5Ec7uCM6chsOlTdDebVVHiv
ZrrxKWpqRw6WmQCThvI59gtG3VTOqQsLo/yvcxmksqeDndHUDQcD393ULQt3TlteK31hRglLAmOB
u6PzeSpmyHmI25Fek9AwGHFca4nolj/OFTW325V5yNTCLCj8UhR8Kh26NQ1TjuDtXiBdjrc6LKyp
QKqJJBWWGQAQgJsYQB3R8O3Mm0rOtVkKz+wZkR5fmtCnUrmqq4TSAP1M1uC3cr+AkW/SXZZUDaxd
HX7S0IazZ99JClx5uUMzpE1NP5hU7Gj0728DC+/hdNOdCjTXNjm4Ikzq+D7f4/s/3C43G96f7+Ce
4t6mg4TWAS00LIgg+xuuu7SJ6SpR4NGivoQIRBfMyHzeSYz4mO0z2WSA2NeKx7kDxtzaE9UzqrjN
3WOcnm4vTO2LuIJtlg9jW22IViki2ZelifHHGl9vqlBy58AK3r+LUbMhrwKJN1z0/73YzQK5v0lH
kswwfvF9NIsLZw/0HQ/qThcLl+tfX6PutJbB2VzKOLjGG1ab3ZGXDS0jr/3AjBvaFonUgSFlHz8A
lMrwK//xBmfoKkKMIpxnG/LQUKSSZmfMBJAjXmR9wV4WaJ1EDfSpccG/Jx+Tk+53i4f2Vj+qNSsO
iAFe4cJ2qssDVxDjA144lQY2Kjv1gUIvdrsayPbBu3hD9rc6jPJbl5Y9YkH37faftOecAQqThaev
jL6Vo0Eai3wJJAY6ZsnURcUpTIgSeV93+aG/D4s00LC5gHDahwXXnI7xuUL6enYcTBKQ/ayIkfIN
yPZbUneD6yrt1TYtVYEMgR+I2aOpF5qTUWk7uD+BVK6H6ay7Xu4hmpIPpGyuvq4IiPp8WySvnI5u
C2Ynin1opRCegvJy+C5GqVqOaEAHmZ+gyJIeZxVm2bXAF8SGFojTG1by7QPnfiewCVZewi06g/pK
p3KwOJXogqCEBFPBF08013z8orXRIlY8bTqdw/+6V9YTxfZoXxd64CqUcXfsya7v5kLBi3hD03Pj
y0SjW/ZlorHFr2UPoP6AvOmZypILpQTu6FCZeyOkgT5PM5p9kpj9z3VEj++3zSDdSSbNt+bfPy1j
wDgD98pVD6kDdM+B66/oS8uF96fKxzXS0n9+zOUBqpH3UImkjdh5OaKYU8JGgo0GjPE0Q0VPKlRD
EtBVLyZdhmUQidYDglpjdX/rpSPrLMAX8pkDEMUPthJagkg5or/7BWjVf86F6sv+cGHCdncdY0qY
adUYvn+CEicQjP3uGDefG72YfYGGDIKGRX4kwcGdsXDrUyrCytGi2AyeJsFVv23lVsEFuqQTg/am
xj/mlEBODRu+CPH20AnUc4JxfW7eiTBoWuyZXAf7W58AGdO0jePY512JCBrQ5pljhsoq/1j2bbcs
k0F1WJ1aV5NKMnld9cDxAz3MmE7MC3Reh6YSua4GX74TThatQBgahth7FmKoscOD4UBzsFAbqaCd
+cMFoy8ITT64ji3/f+Y4Mk5ZB38tQpNYoqxCWcjPuv9SimVGrnj2BAONzCUUuoQDuUQrmTum8X+E
Rg0nwWATTPlBfRUso+3sauSPwYtpK1aH5yrFJc9VM4OVw31YeWHtbc9tpNEjJwjH4sWw/VHb2P6A
jgn6wlG09sbNVIoNypOFNMxDiI84qQS2D6L9eqnDjsw9YqepJosGPVDEePjDGFsLiZVAR4o/bZKC
y1lSCF2nSKWLJlGZSula3t0FU4HOpjBd6S4hzUZiERghMBDYaZjeF7C2e+9y82vPh7MG8wDIU2O/
B3QWrzP449JoG38VrGlFqYrwSLpJdXe8qZ/A21yPu3TMKKUf9G19OmiuNiOZwCf9ms0VpyB/6xJr
TQLB9iOEl1jX17TNwv9bANKNcbEkN3tT7g+lTNVGAkSF93IXyUEHkDsQ8YR2Xy8S5sVUFcI244fx
c/r8on01I6fD6s+NGFXF+jGxQHGd3FrksfkNHRjKycdbbvl33Pr6tHeCjnDW82+VaIbIexEcmDwP
DH/VQkA9SZGU9IkTBPJYmk/PDYMDUTVryGHUBv1Pkvx4xbwlPnRffY0TLBvnuf1GvChH5yrg0Mkt
qcJV9nOdnyhXlqvpRrWJE876O2mvxGCRpoTsNlpInWwl8EpafaUMMDyoPY3IItmkh2fQjRjMelfp
906lLw9NPQn01+n5q275HdZ5mBzYKRM8zk414I/E/lZpvzIzFNo5RZ2zsfDfRCsqe50UeBI8f8sQ
dCV9eNSoDuOtGmQ8cm0WH+K16cdvGNvxxxs/QtEyEn47Ouj1U1gsF4ndB7wrcWo0oSf7GpwkCLF4
RsBcLfaKYCZGpv5KQucw6ObXaGmkk+TXrjJUq7tXd9zSrMWTuugBRyVHoJ0lotKFV7gQBt/Bi1Gk
LqabsokfEwtB+64+wI1AMb5ynPQf8hEcHXcIuTkJ7JooQArvGFghH5xr9Wm6i2B6QTg0q3WQy+4T
QqO2ydbxNxHG4kCEKZJSbMf3tbvLd8LFnroTbrXkY3AxoaXkcreeMrfZfKfp5p8MTAce9YnnSKvX
uh1wNtTY0l8vZS2/E0PSnc7t+esbBTWMGwQF/u17Bz6hQXV78rIYRbltWks7EENVx7zB4ZNzRG7j
BLs/PlNcaNtC+AOB0tAP0agdN/QSi6UdkKPJ8WqhM9xKBfxCek72R/MyFmlEq4S+zI1RaWeTBoOj
pRTxfcKTJoqX5mNggNT4UrMWil5GKbXoXzDRlN+ci0MkKNE9hn1+Uz311JVok/8gFCANoZfhzK9B
TwtoU+reBm3pOacd+tvkMb06MQm1awRMInQj1w8EOlTHb/w177kZgq+iS9QNir0Z1HxC80c3GKVh
4zmADP3ZCJ2/1+yfZbEFLzMLHSIxm8+5YxxaW4AAiyKS7mOqsCrHxN/jch9qjs7wB2RkeQqqgiuV
P0NjCVc03C3b9PbgJbbda5khh9MUjRhfb4qypgR7iTu35UXXkHhlCS3Wq6Yq519EgR+vCen+wBSs
lv54BNlxXuy3wpo/bfbCxj100TzOgmSJUXowM32rY0/fSoFa58zyHyTCIb7xnS9BIiMks9V/1ZZt
Q5iBLoV7b+zig44ICpdc3vsuBzxAEOpfuS++uxDsUFR7gqeCs4eYAkIz3MWdeKTLzx9571P2v+T2
2GB5BarmNmKMfmgyVH6V6IDZ/XSPmqNHpFM1Kl6UASxels2mex43k5bYTLczJdxoMevdPoMcNQCb
rORORphStLsXirq1XvxFyF9zWwEFzeZ/PNf84ZSfcIVuz2dV2oAb3CL4HB8VLM0KOsADkFqD18tl
5yOyn0VmQlmPGO+q8zdbaaNms+ZxN+qQ7IWNNd+QM/XCpZAtaMcyhXHbwQZSL+1U082huWZvvTnc
Ehc8Rt7uJnI8K0rgiEls0Ankm3EPbjUCl7IQbAS+72I+rGzE9vekvFHOxpDu5zKINaoQUSU0aAsk
j+HQ+9+gy9jMyJ64FGrx2hH44bsKgz2cHW5yR6X9iVEs51GWiRxDn3ftHz08LB8+XATZuyJvMCpo
pj1MllcSvJqcdlfcT+KfZ5yJFC/G1PkvXzEY9vIzpNxyyEZoOBXbpM2pBatDpFNoXffbmzqKYKSm
zjN8w/1jQsYxs5SIjmJh+KZuud0+Ux0kJChJ8kc1vVT63CgOzARbDzTUK8M4v1EBAKqIrhAg+gfJ
uaiVCXbtrFBVmhfr7vQ3WutxKcSWewtDwzKXZEI3xBrG5ybaEC1V3LX9y5JQh6qIoE5x1i7ictF1
SbDY9O7lXGGUxqtAzs13amqDynJRm/YfTYy/bMLzKdSwGsqSCoe4HsjST9WVt/1mT6d+614Y/wU0
7yhCHK222AYie3zBhPfFNOfYuppVktGyg7KIMJQW9VSr5i8Qake3Pyg1mofie0YDRju5RpJjh8BU
uDwAERm2+JOE0dUd9EUj1fdgMERfcXCEAnggPPwS6qbsrUzNvn06jbYpW1oD6FaalSrYdgXg5BS9
pGxzoscbXf9gjK3dF4mB0PimH0XBy9MtJj6y59Bur8aYOUFJncgDpKblOubF5dcPNbZgoY96bmr2
bjcMTjZeCbVQfH7fy2AsWUJ5ar7csQqaPsS7vxNiQ1zdJXMmRYrtYxVN63g24CVrZPwNj4UA639d
51WT+YtuGnR+KryMZQxOO2X86vYvTcbKvuXvRG4R2XUrkO7nmMUZGRxpqiQ50+OX58ew9tyyeks+
N92OLy2D5tA9KAiqK3ekD+rt6r5h52Ril5I9CDKCnJW2rPPbCXFQHO57EEVKKnhUwvxzPPNlvVs+
ClumJv3cZYWPmdMWqajpiGArhgBRRozEt0GzFcvDLoyb8dec0D/u/YvWcL6HdV4jaTxgct6Aopna
xfmFxh0y7fLA3zaMhVUX7vTyiQUipkVugqDdU617Qv+dLPYBZDpros5/ok1Wi+qSltZxkIo5MfVM
zQuyjQkXqc1Wgp+A8FtHH84Q5AQmNIwHVLwTYJlpS3me4OuYkBaoBd0RfYmOxEjmgkgWK0DHMXhx
nyhdjk+X9LC/cep+PpAAKdO6pAfHMyhz5a1nvOyyc5C5V55Tsvt1RbFutdjPBJIRezkAS2wKT2Cy
PGbqNf+km9CTSqhEe20YHj27a6ULOzY143sWz7W5kg8uXYMeXILgBJRJj8kIpyY+P70Q7TFOAtp4
Fo0Dn2IerPIz1Zi6htOCOkq9UoY8X6IylYQZ/b2GdgQlVBus5y6rXM/+T7mA4/e76cb7X3OGMjuZ
eaprW3phNzoaIgTpj5K+RsmknvDn4nFS9FysdnFBHKHDzHQyj/hSn76Txitqe8RdW27/v5VKxhMZ
WOnA7YWTH2+uerYw9gYxiBPbd1loZqPpY+//Gk92jehVo57Pwu5fKGyUWNRCXOMTT4ytbcyNtmiU
b/i/Cnprk7gazo6b8NPu1c+nwXdt7x121lnpkRrgbgPaQ6oH9+SzTi1y886TxuDe4Fp3krhQow2j
XV8mB8uVvkSeFg4hBQIC1j0hNNcl6MfwDJ7fYcn18vymQ5j18NbzaHgN05LpB9YNcgd4hiQeimRm
tde9Qp3s4s3jLpUhojuWrUXvB4XOoFH7k9cXD/8pE+IhqhmrVHFQXtmdfHwX6mCQ7guY4ntP33kA
Ur9TKw+7oVRikyjVBxR44gFR+WFxvQPGMhMqUSp+rgLTGGBeJfRfwcEJZ+r2G/ZrEyTT4OyShGvz
vRREvsSgyH+B/ND5wQ1Za7Wi2Oxe57nkWSG/El+HxQtVLlaWJD3P6kMsg3V38X9Nr1JBNxaebFbw
rqwU2Ckf+tgrShtN9xEe+mnUCsRSRht9XvntkJ5usYO2mYC2RVIeCoVKyUjNS1+YuVJRac9esdZq
jeGvk9fCmddd6zllRcyXMyqb4/+XWU1U4xvMMz9PuXOT2DxnufckgyU3RJfWfWV41J0B444riEF2
1vpYpr98buJF6J65QKmiCYqBndaVlmSPTdYH9YAWXI96C+I0ddqdN/yZgxSONsJYTRzaeIiyWHvd
L0Be3TtS2K5JRx2Ft2ht4SfNw6cTT9FklNKqRNdRi6XtNPAoTBkRPrSp0hcoyq9XFtC4+S48ipsT
ULeoUALffMvcVcvO2SV8ERTBGloPYaceGa5dwnBgrWDn1t8GRhLXo8s6bcsn4Xnrl4ziNMIsdblm
XCkBU3u1kG5JFSDOQzx/hGQp/973u/aKuWx+WdOm+uKTMcYayXENDigntkVm4LZnBkNvxeug/tEk
S2WOPoXk5s+J9U6m86voXnoFJakxXidqrl/7nKlJ28NR//S3jkaBX3WpIehkw/HAbLaEIwDJpz+t
YKDfS7PUkcQc2LjGMJTbWsKL/aE0mAYBOYnWpakKikTQe97vOPB5KC9yLugFstgIMa7XzDdWVqO9
pFQYenyclCjQSsMR7YXf9DxYSjS2Czd+3r8l7QniANsfrGgAqIn09cP++HXz8g38KnVjja6BmjV/
0gTXUI/LwauBoI45Q0Ws7+FWFJqoFfZGl2kETxLRweBBW63bSpuFA/hBMzq6wFBTLO+ZWRsMrr2b
WJGJIyHGqnw6E/WuiE++m/cFTkx2I0ndJCWpwu/MAPrea4POqlplmKlbwqhSzSro3kxipajAoIDa
woDg4czUfvRkiB72m7XRFzPtv+Qovxe7DMvnfOc93qt0NVjURQSiNtTdr1eOgzGXBE0fdaVfe2Y9
5/7sxq2nymDx9gJa+MST6FBsKSpUc2q0QFffP9G9wGMo/mVBQUa1c7/Y08U/A47NgqHGD86P497L
ZCkR1bjWx1XwErMETAyaWH8XQ6YPVi5HysC8+wlwMPrnA9aHTUcKD6sIg7VlQfNuh2Nv3i7YWdkh
rjmFwlt01xDLj3XdjgHVM3gnBc00w1pWO9grfAf79zjId2H1ParVMiCDnzrrZrv83AJEc5uP4/te
Kq4o2Ky6fyM+cX1GchuVAlDSrJHufPgKm8Z8aNvFuDoXso/myMpYcOQ6zvqnr6T+T+SIJQJNxTvH
hi4gPmGxUwQMMFicNqk6Qc3CT3471tcf5JuPZsVaJsZ5SSavS73FLoDrukcbtTMugqfTwNLEJQwW
BGPhKuy7t3cfKxs7JtMal75q8NE3Ka5G/EfOpqIEF7IHh/KFPjJXGX/KO6gwqNz6WmaiD649rfGQ
30newKrx0mOxWekvB720MECy1ORR3oMdF0SHzadZ7+yyYRpY1p49zGCcYTa+dj5kLS4MDaqWIq+R
aFBdeaSsFvVt82Dppu+02aieBMaLnxA144QZzDVLXIc1bft8vHSHEYUP+ul23wbfGGvn9uVCb3OB
GRwQl131fLYQaWROXhh7OnArDNF2+RTHoOiHXAIOiry5N21eVlrBvBMQXGw7Vz0+R2VUSMvkXWJ9
djC0Qfhw0UAZEJnsAi9DMWm3O4uT/tduTINCkJW2YSN+8DUuln1ZFpkcAplgOtmmiEBQsxvNEejz
4zxZ8QVtZ/qbeRnZSBqKZUpFJK6pbPFRisYMd5/smLgQOpahKklAJt2IZ8PdUhKBIz5H2EAM1tHj
AY7YPaL+vTfLYdrh+t1W4QFJXO6Vw3SLz7ub0EqNkmKNg6Ecn0OZlmcdIFfvnX+a+r7bG1txj0aO
x4+Z1J3qd69ljut/1k1WUWs7j5I/1KeQzpPcOqtvXlK11GYgAYJMk+/CzsLfD0t0ZO0dMmW90CIg
Ic9dhNUUvpwMhkAqQwJ5/MONEe4zS0SsFmRBqxp3og0hrdAgdfTmlxTuqxQyqPpgSRe2S5QYYZI7
GlKD52Rl26rMxYRNP6JZtcgNhSHavDfe/UDJ1OKavSdqqb2mnb4ASS1fUGFp7PoNgWuCZ9H0hrDO
CeA8tsGYYa1EKcuzsG6wUvWqGesaZzDv466RiK+pO6mOgwx24zxcrt1/Dxz/mK+Q6SDKAht8v996
SLWd+39e2JmIyF625/hEsn1c/kIkve1UPRga+eqoEexKMcciMEyf7kLwXfBmU8ef8kM6CVDR/6BT
4UV1Wco9qZfiKTAmiDQYSBifvRT9pwthlJ3t1H8SOLAOSDlZhBs/t73HEIuWP6jlnAx2b0AjPMFr
oPm+p+GHFYj8KYU744WLSFpxydZnZHwqjNGIlQ+hEXLxmAZkuml1ccQiVWii6dRU91Fg3n1qgwoS
k/IWReTRzn7CFSQ2Cg2jhL84siZJM3GE1gD5SaYXh4wrjQymO9HQg7oM6V3GV1UzRVo+YerL1KAd
6piZR7zlTehSWxtAfs6oK5XuYevHoA2pdDrSduM98pW+cRAUYk80KeiSQs6tuoghHYY3m1zldfuF
Y2iUO6qyZ4/409sh885E/BGWojQKVpo6iUA77YPd+ZTGcRiqBSz2tRm5XZGgpY7LzE1MEyBSP1jL
j0ndrECEvxacm8nILEDLuKsZxYFi9Iz860SFxvbKyeMlXsXR518qrXCBcT4kMnBWxgszH4QQZvBp
YNByje6waRKt9JmxRV9lh6lMUkBTmAp1E3pzIJoCxCI1JtkbQbbpqwr/nmzIteKO0n8JgR5TsMqA
x6oQceBjN+llIeRCJ5AajEfj1pZAxAShtqFoczOIfUKX5ei6Un5zBGKoahipYG9Wm6yxfRCDN7ie
2fu5jG3XDVr1Pnu1U8cNczzU0yTa05nX0rQwCFrsfWYVbC8VGLWUn0M0Qe9Et72JwbsXyVJqSKqz
4GlMv9DX3sLNfBtnTXmPTSju3x34+3clHgLORm7bMTTh26ldQHsUr/uVnaAV8Yp9raTyzb10DPQ6
WrBeH/WCCFLqAvO7cERk+pAEwS5CnZ5LHTc97UJrrqjEW59uzqGc6wdvj6R2+ip8AlrkO1uYxqHL
5r1VYcnyezlqKSDfFQ7/IVY0HicBhE7O05TxooXveBuz8uQixTD94orsGrzrSg9dPBzaBuq1U16F
i/ua9mEiQ6E40kBUFQrhn2Jvjqs0LTLCD0ZLNwwNnJogI5sNhIZTYVZK3e/rxoHe6PKfd3GWrkIR
Mk60FQiyIKcwcG3kVx8mnLFn4LtI00RFn7ZIm+5PMJVH74H6tyDybhXGnXMDyjwqZmKu6tY/ug3v
F+qB5Mnwgzfj81Rgt4Y+EEtc65cPM82sqlQ13TszHiBpsI6Donsy6SesslZbvPt8+mZuKBshdWjM
p7xElnQhJG6d9DmRWLm+8JNFF35i+HmyoFhzYpvipZdMnGfnjYsx2gtoPKr1qh1t8Cyxeguj9tIL
0LzE+niMsASTM/3kuxWUQVIkmugWHbNiX4tl/S+dlRqp6LG9RfYH9agTO/TzehRNNSkrOxZLq2F1
/D+PbXcZ84EHSbSVeGGJiIfjizwrzfkSXsTwubjszYR+MpfittYNwm3keBMIP0DOM1DkDA89A1SH
URQUY9h4Qo1IXhX0pHqv//PmdslazCANdaPs1MKNoF62BlrEQU0EYrKnPWXaUAu20DF786/S5f7M
WdK88xkk9ACsHpbaCDeArdKPqo1xd+cRkdD09hbn3OyY9146RFo6FgwfoRCN2KfwEPuQ8lTWaJ3J
Ax82w/XZFeWqluCMUbixcFk7f6Rs6+pvQrF6EbEr8LKQyxxcfG5M5wJuQ4DmbL9+2rrbiCcMjV1k
WtWLW7fPOe7rpB1Bz9MXh1p4ha2LUMREbCFyi/4lmREHrRFZctf8L4H89O76MiepMwNchmPchsev
VHxqrK7wA8FI8FJmfNiPi6e/Qhcm1mj6RfQcT6+PRcBwqLzv9YCfFNvYin5xgdyc2m5liin4ikyh
+dWdoqu7oJSoyl9qzTeImJb/h5Akgkzts2fJeJErBo/XyqCc5HNtgO5qUsMX3wSQSTZbJPJZwYSb
9JHNwAz2EyL5Gwg1TmmEFRlYSJAXm5vL+ekFetLkL0ogzfQkAODPgXf8iiuMUagEbDKMStQeZhsU
7ibfRK03w3MeS5dONsc7jyidBfPxirGwgdHu+bBsXoOudkSUyt+4ne4MnTwXBADJq1TU74QUCJCw
WovAS4CnBfVHQrk+uOY4eX2zMtDI50B6fpqjG44vZcwpDMMzDy/3IX8eWrvv4xmHH682+tfgkb8y
q3MHDVLvqlP9vhAgyP38NgJqbB8mOoaR978gFPvTetWVU1dRr/4R+1DrnsgTaIL8pzHTMuVoDD8X
Gt6kFgXUJ7p6axmSoR21oGH5+dtW4DrAjm6pEqXEQO0B9K1feA4o9UP0YaPjATE4T14sPCnWYWut
/GzDIhQ9Uw3wUkvE/EIsmhobpQiWDz7SS14Nv8HqJwVWSRlEnEHGTSzr9zsu71r/PntZTw9KhVRn
vxvLH9XXDUL6k6xOwT6GEb4gGHD9R3tF7yeoteEX1YW42/4YCtAaTemGCUKsIs0AHasM4dgQXpIE
+Q4AZe16gQjuPENBNG0m9TzpAlGy8/mSuTkn6tu66mm1gine97EzSl26vkPUfkje3U9iJwUQeBoN
RvjgPMfu++wE7lQMKOTVO9Fn97swSW2UJ0zwy4xjBGnVNlgffzpKJzqkzg6x8g1kzNq/U27kkzZS
mU3GhoEOQAPuVJqPzx4Se9zgTFpzfR1s541f3wxKfMl2NyFzCkZhxSxTUU+caFwovJYocevRvg3Z
7UknvJPUnJUayMqxTvSkt2OJpLWS9vT3hQOeDltvwut9JbKUXcp5hxwjEOgoqfsnaX9thpwOZGbY
EfJ9SKIXEFv6r2h+/VtoKfjzeLY3BmW7y4U0A892W44YKgb6zb1S3Q0GX/Tuc0SidK9Gb5G1CnQB
xkyUZRSimt7AxGhtgFgASkGSBCjOj6rZ+3o4VVqSHnfepMIGOpJHBmygEmRcjJ9rBxDR0/D6dcKI
SnCBQMDp69qERaRMneJdKfQXzOIQtoUpLvrQyANknNkSskFtkvBQgSSkFlvnoCrCaQ0oHIva24HD
p85NLI1+UwBPNiCoLkL2+oX6HiXnDgfNpOnsDcrPyWyUVHRAYsQaUfU1AuT4SkptfzyLopW67kld
NKJn7UFreCH8d8IFXsu22QnUXdQUvpKze0uG0s1FCtYimosf0oJZ+nBUgGVeJGCUo5dAW/DT/eMW
6QQaUzjCHwWeIonbNWT4nYI7piv4TO1VmkzlxGg2dt0QgKpZITXox+LkrdF2PfBhjQBNhF3sw2cO
vut42VAzIJUB7RLB8Bujln9B+FAFGRAkYXqgWrf4NylazYyMKCBoAyocC8sQ5kvNz1JizzfuWQSH
tpkNZUJOykMBQSiKRVS3dDe3Ov/PkQ5zLaWBD0rBZHv0ghvbaw36AL6/oDjMaWeqwdvZq4m3sPO+
oSUZDZxbmVL67E8lATldxWyodp4qIdVRmJOEMhoIYb/qSM8xUnrsIcUvd7LmqNLb6QlhhaGL1Wbx
4Lz37t6BIwJNG3H4pA76JE5ufeWwPEAxMAH+JmZ4c/5gwRKQ4rf7+N1306CtxEUlBWmRSznJ/GDd
wmoAM++bGEbUvfb08HYTjzpSEi9V8FMXCw0I47aEVS2/SJKh0NDk1HvsYExCN8nqXwVznDre1sEn
eLr/PIHQpVPspkguSBVd/W1/Cd0Pud0E9Ughcb7NiKJcZoX2l+tFOMSDP3QNiJaI5oZQ0IxwXNmU
sHSoJrydmdyBq+0N+GX5Dz0pdPKJg3A1SoyKCgWsHvCLDSq83IBMXjS/lRevT7B8O/NsJrOgKSfD
FaiMLOhAoO9vVwhjoD6b6RlLgv78SbHcLuobsrAvG5BKHLpoNfoDBzoN/NB1kn2/4vMYK6C0covr
ioOR0+PG/yj+dth7uxa/Asv22QUMsHYuncYq9YUAPOt41Iy47zxLySYGl2hcBbM+zVqwNxaKA/jW
Mrt9S/QPzdsqkpe7Y8KQyIRq8n3hl/UuxnB4h+xE4VEe1tsFwMJUgRZsBTMFKKP+eZO1w7FcyIf0
emhbByjfAuekdAqdPlLhLi+2vN4NDvUZnLqU4rBLlGXx0lfLLDbJkcCuA6m0v9X2O4WlHRb1D0d2
4wFk8WPx/x+l6UCfp6oGlPotdBHUj3EljDrQtTeFMPj59Vqf9OJK8dF1teKvlEJMt0pPTBZM1oAt
85ZFOpGwRP6N4eh/ps91NeiKyD43M4QuCGG2Lx1EHL5wkfdEH/rCqXr/MI87TyM8Lom+urGZT+sD
t127D2cBlEsFcMtvZBlZDcCGKJhO2puErTh8DNJyxRGjnlpKMVsOL4e6H5AhgIF8WE5R4ZB0BP04
89fDd68gMd8Fy52TZH5UwMX+NdEBrQaWvj2Y2Bktud3tgmVLYMkQbKh7FZd/znEqH/eD3iDeA9jb
DpFHvJRQ1Go80pLe8Lbj4y0iQ2A50TLp2N/kXNZuckW6LnKuq9WHPWlxs3/BrAb+VfwPXJG7NkYB
37annd8fHEAfitZwdzQd8c277THRKdiFiqhVjC9eTn3O0raDV4+mlr5oeHO3VbFW/hgvX3DsyApU
EJdWi5doOIt/aWe+IhqPT9yYR7UHP3FlKLjCz13T8AE7sHYFHUthSKiJTdTA9knvwG6ist27Kq1Z
dBAmr8vyUUj2B/tYMAkdkCqWJSW+CTCTQ7DxHwg1YQiIZ00F4C/DB/gVANfQdAlCKEGA7Y4x9gd8
h+0dqC8U2sF85PS25dc8nJ1aKqBtxVk2dpmBqZHz/OoExRIhPyYlITIatBcVV4rsESVi5Bz4qKB+
WbqdPIHx7kgR3io1PkTV5F/7S4z7ulMnyN4qWmQ3UFnZdIVZfGAaQRcSfEbziThy8TSNYKignutP
P7+McTXF+f2lDbP28Gptr5jaCdVL2qnhKeuHhjugJh3eisJvg5Bh34ey+5Sq5uMDKQRDblJ2/vAn
vvCz7YH6tY+d4VrFK4jhikq7E3k/W60MGUPieoHd8Wi5HtOjhrxhWFmbsrt3DHOVPz8OzrW26dne
72+na3RQzekDuUExx6iddc6SFWtCbuNKN5QIJ5pHeJfhoEgSiOqA3dyggiZKrMt1TghK1URxGXRS
6vlTCnroFsWnjgXZv1gCbqp9FxZHuauSoaoCn8HE27LlmJ+cOBZaabK5eQjLpHOo009QrEeXJEaD
75pvyjzb6MtcysShGjE9Mhc5FFC3Vq9S0OKNWQQLkJbSMw2UGUe9bOLuf2udXyr9nqIygwscEikr
6lnkaoVKYMW8Speb7ejJ7TKgHDlfzRCrBKrXJJNSK9Z4T41aQBl72RUh5SUI5j7IQpeXuOEpVWY1
EJgrakW44pi5kFBQOIV5CEdIYyxnsnCjIPQLrO7dnDkU6xR3JeXorvHvpXWHhQa9LsVJjOxVIJ1T
NElQ7+H5YnldsaOfTAeZjC6DLys4cLJTJL0H2L5PkLP8xmFZlQhU1OCUJqbPWaxv/1mEDXfgo5HV
B639T33aiW5+dAcOWnt+FcnZGZED2Nyt0O2Xyeo1eMoCQLJSd8Wod9fPnbdKE6v+jLRtnkx/wNwS
fCieyIiRyFdBAYjPbkgcVT68Bk/m0SzpfBQq09Zfxj29rqAFZ8x00yxE64B0oKxMExW6At74mKGD
i7O1iyDVdyZl6Jg7/0EotL9TXpnu1eEIxsN6U0eKnJ87uG2Z7eZbHtpdZIkxCwZ8Ap9IAtwKluAC
cBhW0oM43xQN8bGyeX8SY7PWpBkJJ5yTGuiCnF/xYxKbcvfIVn8a8EArH4lxC6WxEG2nh/d3Fclz
ViUFiazwvLdy+wZmjhGx4j2Dji+5ynDT7LprgoQHWYqxTYok6Zq2L03MRziHbPDCs3sA/2GYbWu1
x/kBIoz+AaTFdkw4qUppcfMhkX0gzuGpGk98MjDxNAmCQSedZFRAfgQJ+Sv7FBrb+oc1zbw6sm9A
ap+Xe1Vzd31OiWaMLL+DYm/FRGiZ8RN1F00NwFH3NqUZZ7HQ6tKjNB4PtMbFee9rc/BLRaFsIyhR
EDTSP2h4Sfm8PJTja0AVpnFVKFB52ncfI/B+ObUCXpielEXjKhrCNeNmUcEYML5ST3e8TqLhQxg8
fOkFrciO6USfLLvljLeRl6Bm/MOcIA5izriLGDfB8FmvJ9k2AdHdSF5anQWgyjy+v63Vt0MS4fWx
kl+VjAZRgzAMmR1WJIVt0EfUh/xB5/pNEdfrCA9//1HQnRpRHKaH8acFxCq4aVt7GwfAdU56I2Rs
RLE4q1sOSEcYuGROpDUD0wHrT6HbKra1RjhAyi1G4sjWgHyry1XRD18+EVMm6GmdsR6H1ZwNsWEo
CiNQm+1gWpdMdHorFnrddELfxg4KB2MafJhb6KgxG3IbLpLhx+ji+MCFVMbb/L/nrZh0WfMWBTMx
AkLksG46uwXqB5OI56mwVVsTYxoVhYsGM358Edl3LY9el+BCV+BDW4oQ8+gntYLKCFVfG9/tegl6
NZliha/DFYHqsS5fIxH/CMws4s32sh3l3kuxCGl/4mHJSeOfvaqVGSWG5YKMtCDU+xkNYOUXp5uB
YEZ3BUsAuGXVmQYfO8HhQm7WdIB1rw46nQY6fSnW0sWTJPmJgUWoCW1P4fo+Iksenjl8M+KvP57u
X5gMj1OyzMul/PGPnhaYrjICZVejcpWgG/SgEMLZV97T88+KnGyT5XiEfH4XNPWX26FbWeyWVQWQ
NNTQ5b6ceE6u7GvbeTYOw63s/qkKOJxD/NycIb7DlskZjEtRudf9LqkaqvnNSBWYBfP/pX3ic71V
oAUpmTsflLY7JmXYjLM5A9SiZ7s/0Wgw0atNJUXWgVWXoRBSW+mUYMkwdy3N3ZWKHUox5Vn2F1E1
oar6GCq9n5Kw+GUwoeX2/uA/bLJyJpjoH/PmPLR+6sJcMZrBdBswpZa5pulFgO8K8Spc7mCbb4T0
+NB4h/nhTgUubKGuYYTs40m30Wo7ay5OShEsmz16OeKNLqtQ/01HPqD/hCK5m1Af85w1OcIjgmFD
l4zPQ4D70u7WLwCTvrtyGWTHmRA54fO3k/nr8xcceGxNx3rsx9nGgaQJm93EOGv6be+FXkweNnV5
r/KZwKvtDlU2yvdmAZAxiZ00RdN5R5X6zdHq2WVwCKxYUFWLzfOAJ4FetM99ClnzNf5qPIkaNBCY
Z/jmgK8p5sPf95BVdFWrsgfnSp7+DLHbavp373HSznLot2HOOIdlDWCBzYgvDHlCcW3Op9bCSNe+
DOc3CAWNrx60yz9pTN6S/6+XjfH4RciIPogoE321mG8L00WzHjdCz1Zt2gzPKOM8rL89yCAuVO0o
BZlFimTc6ePtrARMI6SkSCwxQet6hoyn0SEq4KwjlJmnDh31CremrTongFZ3tgiCIITwt5w80TU1
LglcQKMaRv45/Y7Tlo7s3un2XMDtRKM2snSGvWNQNAlgLrSYvzHcP8ArPCZglaY57UG1F5++cCS5
d/r/KKKlWDCOIf3Jo8VG2tB/8gQGx5V1TvnZKE4ln8IokQflGe+w2SC7pdVWNVsOCdlpetcjCgzL
KziLwRmSSQD6PqJ09rKTjbI8uC+FEpJMK4mfCGdVYbqGz/gbCj+ogzIkfKXtqNuN7CrTtOQo2LiJ
+tvrl4b5Dr3pIOY0ByhxgCKchxz0DEjVC2ijy21Y9yoEJoNIQlPxYcxewcVyIxJGBaPaOrv7LkNC
eRO9hUeh9RbF9THqEbUNislhvYMbwX8Midr2owBJLF05T+Ibu1cjzOQ1r3MxaSyBiqCxSCygqzqB
1aB/REPv2+V9qx8oKbhPKb0Eb331fFC4pt/AH0NOZopUZbHnSRaRmuHqbHMR8/5wNunj3dtLj3Hc
3LBlih6J6dqsItH63fAtPzTApcD04AvukqyuX6GyB1wvOgMUddNDW2h+UOXJe5E+EF12PDB4NyCu
OdxiDtgGS3ci/BVqg2VQKBV3jpqqAr3+d5oTVFaBwb8JEMOXCXDUcvb4Z7OwSzOZoGg5Pl4aKNr4
nATbEYCW06ZpvshdzwQYMaMGSqjkRvXH1E2w1MKTBD8t6f9Vakr0/P6ACmW9BKDkh4fwgW9vb8on
ol9eHynZm4ZN/XlPFXr0EQCPsjoociJwKBZi4BPKX91EPpc1HMDXM6SlBQ1URkHywTmxhLITZOwG
VWNOP7SdT8zTg5CNKUHXaR0/RdMCM6y+mTydLB77veIpxxf6bfceYMB+gSk5AlGAO5VJoS1IHOSs
o1KYPNAEvyTb1gAL7XNR5t+Wn/rHqzjF1kX5p33Jnji/1U7VfMm45zJv+g1laUCctQV6herlcUec
ZiWPnGUkmhgO09WTL+Wv4Tdt5/Q7rdi9ZCs9wbKSJgyeE/ebrsO7+do4KSRymIglpwYv2/aCAIA4
H4x+rumNgSOED4AvAO0Ph2vPJpEr2yOJ6uLmL037L39YoIW2twoYOG9NWgqju60W8Dt8LYGs/7DA
oYIGTA+tl9BEpgT5mlK+8hWBwnHe8Dt47TnuhtLrSyfMc1fYqW+IDP0VaRcwfYPLAKbRFBtMJUvZ
0AQl8AbwQozKHa7b2fLlf4Ta1X0gs82mRrdNFuZlomjOa/WYb5K1Z35I6TluH4kjptXtFxGovLmI
8tyjZxahkZErNmAAc6zhWmJJ8P4WhlvhHBhwjeCrS/61D3ibOcprX+HMWKmM9ZqPDd3hBqUaU53U
bvhCILSki/Uz7fKJMZp8krIGUpIeB/X0QbSF6fQBZIDmtKxX//hq1W7pgLeSpvhnwxe7PLW/Cm58
7yd78hgf3STu/oQX3bgsCA3zbOIWdlq4RJFikI3P9fWWeptfMYT3bqGWrreaYBUkQiAlgi9C4DyS
pMfj3GcU/f5JGi1tyiauBSUIibc+QpHeSsDL9klzN/SEM4TcQEPzwdUwA9Cs3xcDDCIQPrznuj1M
wYTEnVjXUsb43gu8hpheTSm1bPQoQSTq8C92eS5fFqP3g/Q1e+sAd3e0Nt7IyECIgdipzFgfrfZq
XdK8+xCelPdeXMsZXVRqpgOU0h8dbVyqDoDOGBsPOid+fgJmFEqpjD6acTndUBslW3dMZVoHpUKo
TYs2OxGNXbfBQmV7XxQkL/8/x7oVKTHkXAXEjSk2/sGJyJXP8ciznijjfoyxoAiRZ4tuag+yFU2R
IkUJ2h3kktirMyBBNPJr3iMV6TTZ82sB27Xd3ZNccbpK7jFNb0d+JENi9prGjVbGfdxWMwXK3YTK
FkpwfF37SfeWvQ7R9c/rCSaJ+C7EWFS+hlSuGDUInQx8eP2JAP09AykjJ8f59SHbedoSMt1HrxN2
bEVXWmFAX6pQwPbDqJMo1maOs//z0u272R9OxPJdf7BlRa5ZKNLG7Tf0cugqiQUVF3YY7e8RloCl
gwGabcQbEOJDr022NZrfNTPD8cDFNIuYTIMnGP01k6tFrjAIg6CimdFX7awVVXHrzhehPiX/NNfY
rVIvVA9LpPMtp02HSFFDNymWIpCzTFS/hgqEwzYYWI5knYrj+53I5Je9j4ku/Bk36qP+eVv4I6Y8
FR2e6wh3jF55fdSfRFslic/7Br5hTVXqgOLy6Q+keG52vN9e75rtOkTUKyxhiSUY+ny+1Tl/cqnB
8XlZYuGb91eJYnfIstslJwezlJUBjZ2BB3mHZKxpN5wDQN48cRTKjE3q9eYDHFybs3iAZF2zbrBA
4c+MBKGURZdUHs/JeXesjFXSSBvvAOvmF7Wi11vBgPUgSAAu4tYjawUtC88cdk9aPA6clcByALje
ntvMnoEK5CFBqi2nUmFJWb7odRQjNdDt10GXFpSzEGCJ0Q47iG8RHOjxtPJEJHHBSWsiuLN0j1Tf
Vup7JMIhmMCmYNAicjPq7CJEdSBL1PSD6pkwWd8yDPesgE4pikOlshgRDuaAhhBofC198xxa60iS
wvW4Ksk0KSRhlJ5rcvUQSfVPFoQeBVMFEpiyveByfM6MnwgbloVAYwfcTsBw52Mz4XicWBzg6AiW
8RsuXNACQzAiqWWmNRoTLPPZeDlqi2VUI+zrnllQfeU271U6daSZlfaUdGTRwzsDVYeDGhvhN5QG
7o3mW7S1AoHXLA+5bwFj+Kdt4kizDr6drfdHoKFyXPNt8Gg9keCetGaeB258ZTADQd9gkx02www6
LLj5Wv3bo6PXKIBhSIBUniBCJ7IMo2ao16maLEBiqTVRMbcydfGcxO5AycwPOyEiuG+PX2TFnta6
p+XeCnwWRLNph32nuxhz5alMzFrarTBB+OgXEqf17D+3keWysJtinw+fptS3uZgtG81jfOOaA0r3
wmzBTHNCyv15V6RR8K6xYcICrZ7pSLX3mi2AcGAWVjr74/R6OXwYGODAMsgD6KohUUvbxxLenRkg
fF4LNjpY3UySfH31D343QkI+Z/E+9CeBRUNah7a+g05bixtHxeTIS5Ys3tbXYQ6QelGaTgVvKB9C
LCzx6UKwneRjHzwx1p/RPpgV/3+TFs50bshVbBOQ3KIyPHn4IiQecGao4Nujsox4MwJDZhOQk2VI
UOCeCw8+wZ6YPwkz7OOAmQW6XuSQsTA0sq906TY7NVzbIDh7FzH7MlmAmyGdmsR3wQzsyoCiA/kT
Wq9ymYkdt8rKH8wpvxyDXmghnRYkPBFGszZ5LYKe9h+RnF4oSLlL80ng0D5hvTUW78O8Xjm+o+Cr
tb1xw6GKxbnA44Up9DNamnFwuHgbT7tqxnl2sAy5q0W67D+G4xKtHSnv6kYVufGVqYU33KtRf5yg
Xj6bwWmM2tQ/vTUs6tAHw2iM5E2yjwiYVZVev9iQj+JA+EoBZKIyNEZ+/DCwB+mtjRrqGgq22O6k
7KCijRzp7S7GxJ+TytGD7s9GP/fomB5VCinc2un+6PtiyZdvpJU3y/cuJViukE+GT1oA9SN+Pd/8
AFmOeBtORqRxFZ9heNoKPgk6Fwj9l1280PZFlgZVxLX+ZqVK0H0bOTTSKZ79VwofllMdxTMA+hJF
zRqA7MXkzooFa5SjO3acSibFl5AtOqPitGryUB1nJA4VnAbkeYPmTxBjsxNRUQeZ2d8YmKfiekPO
D/vljrqXWXQao2rtWXPgZ/ItxD31wMicwb4otl1FpmlM2ycAyvPg2mcn4JMCViHaz2rXBwB8KzLm
0GaDeX8aO3WoKXEqWW0WURf42Fm0aALCI1WrBVu6LECHwtjOnAveez5YHpyrNBctsy0hKXSmE1nW
dK5zp7bBNVqDFkcMi9y8ZS68u7hse3aohDCFBYiUvGxoilMJCHlsCDZHTNwWIJL4R9c8nmaSbVak
IjyyAr+oufwy83snnfDHStJn53nbGIP5lcbL2l6B15UHDTCh7KumEp/aK8bYalePGKc8wFgwgLOm
SqYW8pjET2qCjnwMRKrgmcy5ucq62MQ9q4+eWa0IdGXOaK94suzDOG8uq0muoljoQluSX2mH+8Lp
piXK3poRM0M4iskUJTbxU1R0cM9SXyQngq0U3OmCW4d8Ok47qw7Pew6ObrE+wHeqRzEg0wIiMKb0
PcpUi35ZjC2EytDwqoqXXGMyZXVON0DjHJAIGV5zZ7QjOazGjhpgWN/p3jtoI13gTCsuKsfPow1/
I7xG30GN0QFK3jygElAa3c3rQ5A6S1i2V2G4Bn23Jot9FE0GMct/WCRkGFj23NsOniz0npJOn5aq
ZMvYzUiDVRNch5Wrq60JvMcBbV3tIHxZP6vNIeYn95/7oxbCodfdT/UjG7buAv1X5o5MAMQ8vplk
blpffzUSjzY2tuJbnZhV6NYAQ4ZfQH8PZvmS19hw1tCwNwvGbEAmXInkCM1i8iBxGL3cKXYcmRay
AkwXr62/0lWpn+xE9DNjuOxXOZ3g+KqhX601ZQEFO5SjM/udEjz9NecMo/K8vmUWNtXbh8YJGDwU
tnanORPXr0autsoJ41FnYhgKW/zbKMBGTNjHscySPgizdCpg1n/KAVR72mSqSXGDiHcpFLwY71tt
wTbcyd6hi6sl51JqrmPJ11WAln6kMEsTdEt/CBxzkbZAl5hGNZ3VBYehrSxQu7w32La6IuzCMeY7
E3n/hL+TaYVjwQufF+IEwo5Zu4CXYjoO57Kvf9p0xEk94HzoN82Fsr11vavFlvDk9gLcJ113x28H
Ghw+IvPoUlYmniaZCD4B+acwJcxSnbJpZlD4R3vCfKJNmJbV5XDV72nifZQRs7ArxY/4bPkRsfal
1dfbTFfZI3U57k67BJ71LXpmeRBojAp8Uw3VLwUf4O5ZpQ+TPAKaGyNAeGgam028I+n+50nPBwM7
2CQ1LYFhhEigrjmEH8s65vYaJ1HG6xgEaJX9pidCFddgpdZbn/lDrkfV9mzRouutEDOgnU+YVBit
L5Jj7a0l6vbjmh8ckVtoooJmHYi/ez9TosYR15WgbksGye0npWSAOHItGLJCSuiULZVr9GEjf0NX
IfOIGo7uY9XIpXrf84IrtQoG0eSY6XCI08kiKYu4rbyB48drIjVslsUAk7fuU/vPc0Y/Jz6bmETr
hDsmg4ebagT1rDkFAXuh5DaK7XysFaj/bkEz80UykHGZ7PQHhujgwtXQJ/z6h9ZYhmJr0eraRzfn
IwJfwKdkV2ye2JFD/x4lxIg3iowloZtYuBpcd3sjN6+VCDZHhd5RLJ3WJTuwebKrwKKuZZZ8QVl3
PICdK9JMnjwlT0znw5ql8hXbIPsJ2z7dFmJvpeEwutYFLfMjuTSehPj0jXKwnnc33HVmideS9oSz
CnhS4LzEIH9CHtZ5om98ZRmzgNwEU4VUefeBS60UG33TBSFcLKlTKYGyW6HuA6PQtUxRb2ul+nZ0
u4rk0Jla05jGOivnkkxDiGV1+Y3SppecY0KgsQzSSW9l3yrK/k43C6VYWJ3kV/br21mGXRzzc4Oc
qdFdVyMPzqbNU/0mL9Q3JNzm4Xf7WJ1t8jfQEOiyCUX2wWiEH4N/SjckNg74D+cmTazVmRZyi6Uq
I7vGXS+4IkYFaNhOxWojA5C1ztDANBmA8f28va8Ain+Wb10tTFKkGZ9LjvDuQgbzO7B6WmWRt88L
zjeliHzUigriQSSjxQ1kAuDaXKVskASCERGEHrVntbWHf84zADOcj3v4V5ZdCcELTHANJIH93n+p
hIaS4WbK8whqFZR1qN1s9bNYSwBL4QIE145hodCXUSUB4ZNG9MsUOrsAmP4ZqAtzNJbxddfhB3uh
F4YAENx3PCMzvbAERh9uMvgqSk3bUO3yQ80A3wr1cgEIo3ksbWII01dk2brLpic5L4Nlnio1EMNU
SVrtPnBkQE3C3RtMea6VXA0i2Wpr9bQ5Np9LM2W67lP/NT5R/LaizwNNZhhZJC77vZ8JKDNOBlz7
y+SZ6dFsJOSR29wdSCeQ6E2t3OaZoEFXyevqfE0l3jiMk81F4Y/k7L3KxT+TjRo3qffj0DSF7PIk
OIlvuDBsmFSuMa7fa91FBsfIMYgBXrFHXDQXNubWjvpu7Ei6J59slwxmfe882lKswsal80gLGsQk
T+7xj73Vwrei8fKiVjBkQeSLVUgB2tB/yzVCrcrE+7fk+Ai2cvpSxvEhoiEF3qlg+NU5CBRttCOs
R17mBiG98RSWpgNNTT0NBa1Ic83HOBaeWpd5sTrpkZbHdFi4SfahgGnBAU6HIxyYEnsv3Bu/X7Em
SlAW+kmsDuHtTK3Yutk7b7IWOyvSYX0Zv2XxmauJWtosiHNwt8nkZt32Sp0UmWhYDnx/wdLMwja+
l3m0E590as7Db1084DbZj6qaGLNQzbouwIf1ve8wxlWMhHI1bxiuLU/WFVKiK8yiQsgqEoBllUAc
EgnHfullPuvs55rhkDnVat+QgDeP1O/VPT+pFVJQqrpZVVQVvWzGsZ0s++QgqooE3PfSKSgDs6if
xWT27iKAk/SesaPN658u4yG6BTlS/REErFVX6mtYcFDKvPFyUBC2+fGTAiwoE7+TwPuBD6RVrUzg
Td65vIEuDbln0Hbpi5biIeYT8WdCAAgJYnc9u/GaJDVS3CEfxCooL5YP8+9AHaJ/C+BS4/8dDtSh
yuBoi2IYba3ji8G7hAtipNntUhP+ZYFokrN5KFDABdPWrYIHbf0euwaUkDgQD2kBMm8951eqVQgM
nU4guMi7bH5xarj3LwDc/JE3AVjGcLcXtsB27dog0yjnZ8u7Wj8UP9Yt4u/8fzg1tCLkuQvJ36OL
v97SP8UImxbMMwuzParRyDmAM9WP4G27tZj/Zfd9NLQbX7XbKkpG26+A9kbxUTsWISZlxr+0aUx9
I3fAo7MD/0/PD2AmPVD2U2G/oh4R8CB2caj4sWMMoSehoG4uh6WajJ6yipEUH5hyYH8kqoEHNKgb
BUEaMjCWbwydG5xegr0heHxEVQoY/IJZfn3oUdaG7kDfLn46o7bIhMAHhYCWR+Sv8CkPNMuTh2sS
jihcJUG+nJcF/sBx3oo0hBTUk3I9atsfqA8FiViCrjIoHw1ZUqV3AwjYNoUOIPiWce03RZJ327Ox
5lNuVNbUQ1DZNkhr/eyWx9UiqxPd7tX8zSCJkTWpsZzjThlKd9Lhdr/yRJ8wAJ5zwnSU1RMeBMMc
0Si54A4ND58hW/mKfxVtAvyd+67wKTjGTZLl8OciU173ABF6FUIGxLCb3w0O9FVgBOGJtoPZEBnu
OiBAiVZiElS0FoVdXcBIy/8BkDdhVMUHmGuulYH+Gm9tmNp0wEoxo2HZtcqU7yPgvmmiyxtUGAkS
Q+7F2H6XnoPRtyfQSP5AOitnJf4Rg88X1EQMWu2ongf7tII49es2fCIUtZneNof+lCLQ5emsHHgd
N5hqN4u9HHtqT73x/fTc+6xbT+SfDdf5uJMIMX//Z6ZYd7GdcLvqZ4kGreG5JlV9X2oUpmM0xI08
mloC6U+tSVzm2ahTEG2sfspiVKjaTwXxBXw7tJVLevPnBpuY1Tr1DKdnK21MSYuLOBjlGIWzNkNj
5SaGgd6mqEk+wvva113yHYOUMrkoIeo9Sv5Pn4GYARKbJU7UAdl5pURFq71BX6H4Yl45yOEcsqBN
QL5ujRJ4MIfipIl+Wxu6KGycA++ywhuEidz2wblkKfRms7h3Eh55uJTJrojvydJ74S5JoVNOkXBl
MNbiCpIuExwwYIqTNhumd19XcwcZkY4jHj5RzPU1L5jxex6IQ4aUf81yKKFkXl8gRkmXT/cAT0OS
Vn8wXmL7VrV4sGQfEcDr+h2bo99g+qt+lSHSfimAafWWeFEQGXm9IIMiAXuYTxAyVYsCHIPzuj3f
komgelYFZpgfim1pj55Z0wpbTsbSp2n0vcvYlBQxnWdsjUA7WvWz48JuWnxwlaBO0dTN1ftWyBHa
jUj/RKDIp2Kok3jKCn4tEYqJOH4996IVhrtT1GA7i/EKcYQHbyt8ghycow6zFg5HEFORPG3hVkYh
DELc1KExYGjzpuw+EyjRBZX7RT2HJ+ESnReOtfn+Yxdt4UWjjAadJkZHlIML7eE2doGjcU8wSkPz
zFSymllBp6nWmm2zCcc5xTRVud2eUgZFihmB1eMWKoKQlVpKhDRfXXWkKPSBMn4pPV8I/fJHOdw8
hT6hn0jzikznaOx6ondJKcD6VZiTu1IVk/v1lxBeSx7ciOcByPuv2XVt83mFq/1awKUSa95DT7zz
9X9HX1teKgZSu8yxUPI6fYfimf+tg4i3/zyyzU+OeRNWzEuD+hk7mpG0Z8PMmD8zxsIUCSw56zRr
MoZN/Xo/ipq96Q3F+QjfLYSHRT+ucEzesCdA8TmVJ5dM9OxCjbptIEN8Mc9AezaapYcqYYQGIw/6
fcBWOzLDXxnqrRLVzMreTwoOfJjbknOdTAZ/Uzm2u2tB1xYJPeCEiMZ/bj/syz15YWW8ZZZFFynq
5dW9Kmseq1dI4Z9I/IyHfzigt/CgQgnxvT1bgzj+mPkF3wqeVgEQnpvfy0ML2WrvNmoGc30hJksJ
1jJGy+U1gWjgZ5l66AFb9AB1zoeTm6OQKkB6tlr8SqEdWcmrTQXVgFU/zU4G1WYlEzrlWsm5y8il
1FUM6v2A/zPVQu+ljr/0K1ZNr6Arrr+Ayib8byts+pxSP9sDNIyzFpE6geVWS6I28GzKlmusg+sO
jVXHIlA+6lyGhvBpkEK3OM9XXqBMXP8N2XUjvgB6+en8IkG0SBqn3+wauGM0GPd5cOJUM2vcaYfk
gMAZL7i2EgE5Vc5meXU3lk0sSqqXHojxA9RFpRj0MUAc6yY+2CxQz/PN326CHX2YACL97zpEdZgf
aq65KI/isBAArIr2VCspIj8fXy5k2S5VyQuEH3F77YaeGTLXct3/NYnqSbUB6rb95+AwNUQULH1B
akyZzWWbX1ph8DXqaryYnx4fAjf0yco9Ni9eoKqV/6B3njVNiFKWRryDTJVdxiwts+2cdaLufFw1
EfF2mkifeMHzwlx3GkG4wLHQFHVe2rNn4XdqHjIU9+/hqa1TEo5EFuihgdQGki+WEta6q56mM6aA
jvqyCFgc6/U/kku4htH6/xjNiMwZsqJVQn/3JAXh8Ce89qH9F29E+3ClYWOEfQOor7J+ySJUKHDH
TpfAwnDD3gVtE4ZGvBK6l83xUw6109ZwMe2pNkpDc915qUhX7GJsqRglUkL7jIsPEK/D0xToCj+G
fErQIsujMIEXAMcPU0OqgOCexz+xR+EJNXY3eLZyi3rmrGgTjRrS7T1qW3TqjB5g0wwbNqdlGyDF
tS0/Yo3dAgngiEKYeUwAbs0PfQxskvlikZaJpBaxN42cVKOxxWpYDMFysvD400S+Wxc3oaDRSTOS
ZJr7Ji4UFFjoZYSDSQGhi9A32wo9nbMwJ2ZVGuMqC+VXqO2Dm4lPiwL1YgMXnN6lPJ2d3VACzrDk
VkAfspySIM2aXQsZBPAsexlUX0lqHlP/n3KqhUMA7kUthb+7xTKDxQPdTAoDl2CkjtNi8Vsh49VX
05NvCP35amAH+xvzqTHTKxv6Fpvft9rVAFQjMXoaX1tK3Wxg5p8Q9UBNj8iYt9TGSDD/bSrVWfvM
fjPmouLd92DW3rNKoNPxGMExm63VumWDQfO3t3euFVNkIXSl6q/q660eab4pi2Hj6jBAPBO5qZLm
xUvSAEJe74/FmWXv9LI713SouByumFSz1Odb7dc8+MuVbqd1fNp27L2Ef+CCCz2q34/SmhrqJSsM
bjXUG7IxjPcLVa+4JcoabAE2VK3FwEvi+VTTY4tWJpTD+Zl35/j0qj9tcvk2m7PKXukplBumD57w
YnbnLfTRvPi9PBDQlhAmIVjqK3kUF0UT15DBUbyQcfRIToKr36XpGQgWBE5rd+WwloUVl8J+C9O5
F8+LutdIxG3iL28lcc4yAbtyJ47NpG9VhtSbTsA5Qv0WfzIanjE0Gmr93D9dnEepE0LcU9uDLs8u
tPJUPyGHXR5lq9ylTSWR27EzyvINQM72jdwstZ/aw57+8/yZTopN/3N4PO59J203Wjye4mGhyTAI
fzniWUe5LAYFWHyQ8hY8jp9CfT3k6TR8pK1UYtGLZnWg4upuAnetLPqzx2h8IfhVoZu67Rco25jl
Cq4B/m4b7GOh5CE1Xb2Ldz6RSV8cQeYulOdgkAHLdJZ/l1hgPQd2OcZkHlPMSUqseZvtqSICO09X
WenRvBJmbUsJ/jwI4RjQhW0Ia+SS0GHfjekTXhYMmDckECWTQiQmvkBP/o8lNjR45IKQ83Vx43qx
dIpVJIfAJBnh4A4lmKPb7mRh1tMp+8rjBTaIF0aa2DR5oQViLOri02sVjdBJjkDSS9YKqA6IEtjM
6nzFQVmGA3gsFSEUCMr3BIr3K8hTnxPMK1hRYIfTO96Lj1zD14o+M5KP1Zgicbe/MxzAR6QPooOy
lRrXo4kPEIskHetm2TH0xcsEpVH7NCT6qhwU/J9T7xO6HbkjODTfqNNW3nZ6q7JXsq5jaTAZbYfU
ONlI+3kBl+ZLhcNQfOXq8ZH639nhUX1SE0ChEQYOKN8xAknJT7FUh2ILkVEBqgxeB8lCSvHE4Bra
w5a5wqkvCaqgKD62o5nvqzHdUgKiENiblMry35rh+Z04GrPYANjletT/HBD8lnd52IaNZfQciYIY
jsCpkQ0lwbAGQLP9/4ppkEeHuV+volxdCd2/b0d0h+FFlz0f6VG7f95R0jzvPWe80H4OP83taB3F
Ma+TiwOYbLKx/kVNfKwkROQ1g/CAb9BlZD/34AiDmrPV7XuAytUH1hm+YQYUpw9/M5s+Vuv75khX
cXkS2KVdO2zQeDilWrZ3cFVyOHzPc+Jg4bTIofGqQn6cI5tSgo2t4Fx9IBK6P4bak1V31OCpZMDV
I5b0FzWeEqqB3G1H+vHrYj+IVoGsFWj5s12rHUGJxCX8RwAcDKpasW5j6GI15LXxdmVVV431/AtM
iBD8kGy5N3T2FFFVZT0yeRBQzkw1wla+5Jk5tw+XoBqecQY2BfpjYhB9IZDQ09d3l/MyYN9WjQxR
PA9iT1HDvYc4mbKkU/ka2JTpFRnoIWcdLBd2exnHsNnhBgwJJJasR3k3N6z38Pb4D761VbAWTQC+
HlzAKRNFD/qqTxdmWNs3sMWW5L3VF/MMOL1/GJBsvZrCPNDKJJWvps3YLcCc8JNZlYxPZ6+zvlBT
/RXj4bIf748qoQVXPvitViImP1UpHeTlbYpFtPXUk2EgmyYdu8LZwT+Ti9aR7CvNktEGmVwZjAU5
z3Qwk/yETOaVh3Z6wW9NLViaFoiz6ro48RfAFAJ2OSUyuhm0y+FXlISggr0zo3B6Qhi+yP0nEwaz
O/JmscQjV8UaIqMXwFCkxZh/tc35OXOihzACdbryt36X7O7HvOyruOkpCekWrgfAh6Owa9Pru80d
xeYfVyuDP6bQGKHBZ8+2cRZuejf+/VAGtcN5jblu/ge4fks3K57DVg/hwB+8ctLJjrPQPIfChUs6
QoHESSHmsk2XJPmdvpWNx+sc6tIAFMgqbosccIObhftT6H9jtwL0sxHLM/VlNK9rmZXD3wT9zplD
JlSCqXnL3WSZ8Dp2jY6jqgZyxlA/ZppHpZchmX4ysgKQoEZ2qXkIei4Owze50pbG9oCKKrFvu9Jb
DHlKqxw4WQ3cMnBWk1vOf7eAn0kwRZVHpTc1djyGFRS20OM29DH8+yFhnUx8+IhDaSXW+yKa0GSy
Xy+OgvoUsi2YZX4uXcgwFWiJWLW0hH36YQt0cHne59NVLE/4DhJYu7ickXyOt9waa/GG9Gu/Yz8t
FWMZ97YhwiZ6zVI/IL74WnwrGsAKXaI8vz+rXU8YN6Jy740R0ohy0cBnlE7NASjCAugdeODahtLU
BQHPz9A5Traytbr5rcY75vu2o0UR2DccQS3ArMDYS/9Uj6V3plPUQ1a3TOHYaovFN0l/n3N6MfQA
2RHskvQM6I9x7BbkJvGwOLTKgcl55p4juh/Nonw8qRYi4i1GTk1bebBO8j1h5Vj39pVzCKlEIrDN
kEt+SOECApzt+Ya/OL/hJSGB2dD9OoAm1jpc6NLKoj+VUy/AeNHAYVD3G77yZifGKnNFxcl+odvI
aD82CChVWwfg8Q10zeSxR/VVCK8faW3t6WaAXxd3DfBJsYpty0ClgDfe21hfGo8YL22VoRuV9HmU
Z3cxzn5Wg3NRnZz3g3+DQxVQgsTC1q1f+QGFucF6/z2hcHYvo5wKNNGFc2rHCQ/Gktsne1gje29e
jX12c5ItEjkHCk6d+mhNUsKH9knkpohXgEng94tFEfw/Wa00tmKI3YkAym25itKkvl3ynIPGBQAn
31iyH6iuPJ8/5jRp/V8nSTS+o9rhkT0/ri611YueyObAl2AqR5CyfXzaDztHZv8/7HnwNv3p+0ge
fW8FqAaoW+gbDf2rBonpL39aToOpvbTNjzDGrz1mrqmPLOwwwzzBiqJu9a9BYbl69HGYmn2BsA/g
0RZDUdfL6dOwiFs8wHsKl5KZ5hQsnkEgD/asVV58YVfOhVXLk+6C6PAwKXntb6/gPzGzT5BGskuD
/owKfB8aYHqL8NzXJc1TXrnUuK/MIaY3A9K9SmSj3nY/B8H8Xfu9OqECH/Z1Ml4eeZ6gyUmMFWYC
ev5owmOzb1UEQDrGHUQWaz/9ruB5t0DE81doqfzqedzMC36KuIB6gZffvYOtjNas+n2zlWAz1ror
FvNv0kDknBZ5YMgC0DTADXbRQ86wi4IT+AWxaphI9hMoNieiPtdXy97n8Oi4gceijDllf61tNEJq
HmKyB3KMbCWanh0aBYsW434UNvMiZRPE3O+CuRWIF/hGp2x6YcVMz8EIT5KmuO1yMH/nGPpSvbUm
TEFpsE1r0j/33RV7ysu1kgocb225qQIeED6rZE/px8ViBNkHZVbDRLIsAtyMgWrjiQ/1CIiuh89L
wFOubI2/JgsPdkEsqMI6zgSHdkpOL9PZRfBOpHaboSOEhPHnQK7/fQL1hGMHnjoWKotCVKmKYZkS
9Zw+Z2t8hHf4UsENCAUzqnCXx34TLkQudLz+Ve7j95NmBmXhLGaNL9YRcTt0pWrP5Wka+/lozxx1
JajkQjssotUu7D+VFlxiRywO1z3doC9zfUiKVhmz37GDQqe/UyFSLPjYfa8QR8OA1WWt8NYZkAyR
L8gYmBDISwEOPExnq++9WNYHSXC61TlqNvW1XnhiQPU/rPBHW7gL3lIzn7uvmM36CXgxjK2j0Y9v
yz/J/d5hQabhiD8mZHcbiVxA8vfkJBIhl+zNDUiKKqxY6FjemEZX+R/aMQqlBNBk2JRYGU8fKvGM
hnhQjcKfLloxDe8SliQmR+3pU6pxItCzuS8X360Ang0uv+8hfpmMNnWMJVYsJv/LIrKvWjd6rCY3
0sc38UtB9PzVE4gG23sivbC/XBaVlitOToYWLgwrFxnGyiL00r79qMLdagPpMvVoDayJtNIigUmu
VtiqJc4WpfvLhOygPPtL14nExmYijQ1UUSmKkvcRfdCpf0nZt/Tt1MujA9V24rpWb0QQ8bTTtGwo
HtlV0c4DfLPpkwF/QjnMSmnTnT8D0JDB0MHICk3Ti2FF7IOEltGg6KqOemMoir+OqjOFn+U5RUV5
PsUxaMWV4rsfvyJtHgQGMiQ/8z8TAm94yqjPjX3F3htM4Wprn9+P+VN//tlM5DvVzZPKLfKFf+ub
SDhPAexGIarhnCVFyx7bbvgPeWodTHJwaqokGTC6QSwlV7jqxJzGD8/9BnDEdVHwPdESpdPwWQkw
8R8U0qY5KhzOca8I5TYvMTQfYuwWUraTaQmVfPKcW0cfwy8Y1GPrx20/fqpm298lAv104OXJyRiF
8L6sKd/miHSedNigvOgVNAYbm16lAzJdogKPUA87/RqstDRlfcFGZqetz83j+tAeXl2CMrB3pmEx
/TA69WqHRRvJWIEKMrKT2gCbt40qSIIn+YtF0mJOxB09yLqSkGpUrqajYpa5EC7jkspTAJkl2hWv
vXBg4UNvzr3kc/A66GRT7uOOriQ/ZlbnzcAuUzd5Z1Z7MKasAwazXkYVnT8xy97p4TczrqVJQaf+
I85qrm/HEI5NkdWkAnSnD2Qf4EzZlJ6zoW1p1C2YPGAeQ7AeeJ+GcyFDjmiGYuddyzqNTpCNG1+7
hykY/M6aQVZ2chxeYvdkKDB/zjKCqm+b00hP4HxOUspjEZMUddbROM05i/lXshGx1O29PMeKvtyr
HwXdspXGbg8keVAPN00exQKn4zuDouXRyC7spCG8Gt+VpRQKdDZBGDE63hfBj0O9JIcAeHZaSRL7
sT22d/tMRbf/IHMi7CYGQOIuacX807TgJZw1U4gCcHY59iwzxzsNQNWNba6o5HwSroS7dUyTUnSn
OKsy0nyJ35XaMe1e25r3dorw6/c+2QpU9PGWPWiWMfslFFOEx79ebJqiARYpuoZZ5p6DrbIt/RaP
O0JPy+av+eQ31oDPGaY5UugeBsZvseEeBULL9YOgC8vCpingn7txrWwsD4RAx0gmwY+iYQJtSb4h
jNEFXe8NZ/GU+xBbF2UTC3pIg1m6+6EoyI8XTq25b/5W5glq1lL9Q5ggcBLAb/hD1fecraVMRVcP
Z3pyqihhs2xkKvTap9zUbdhITfSt2q1wGlwkEtg5aYfU7ICFwJVibKUcAnThYIfqu6mUdBh+czVV
sk2OIDuRFz6+1c1bhn/SGcVsNROFmbMK3ClvFwCEH73jVYbYAZ8gBFUTCYDl6ffNDeuABAlRsVuP
u/IER3tlPVJqOj381Ujc/WCvyF64M5Z8mv2xrPb9WkVmEehyQbUZdN8a3DFVhEE+ErW6qI+gpzWq
RWUx/RUzNZHEqat0ioMDruyYYjZ2udVcVDkUrBaOlJyNdktwKBRKxuIpuzBZFoLLVzHTFsQWKi0r
fClNjCGRxTTkmNPNE6C8pbku9oBMDz7PsPrw9fifS2SeZ/oX/Hk5b3+rqffxywg8l+uhxrSGXPle
aZjvfvIf9uaxHXxLxVyGKvAdUbfAOare6+iQp4jKkV1afgsY/2tql2pwFcWuCoK6tuG+Rvsvg4By
fafud9y04sbxt04L/9yb0vqMzt/QeQWZxDjB73nSCRx7w3uvNXqqOg01ak3OsOqMjkY2Y1phKgiL
UKTo2Bby3WtK7x8kpea6/OD/Lw7UtivLVAAPnZ1vkMyZpSemkbfz+6wIfoItvKMxz2rkC+QsQPv5
5yx5MDTAWEZPhE9iKZYUQhUvhL/m2wAsCjyBdhOiKuX57kVJicOzNU171gDYJoZH/HbbdR46i2Lp
zgy0ROzrktrgcxpen8ynOXfxOC5Gu0n5IWOOY15avzizZ04bLYP/V77uG+l5kLlFdWlr1H2ODQtN
+76DQZVOaF/Slfoo3FC7WAaXpR9WfH7aCF85q0Ed7GSzchYgiVbx6qMG5ghQHFpW4mSjqgcWoWJX
1tTMaoP7TdDCJ5Kfypd5J05wwQjKEVuoFXSSBMuNOdpGNrgJhoD/m6qEZHM4rUijPLns4Jjv3aKt
CyLwNzH+SakQCeeucngA4u+iZbULM5cHtd/EvncUdpvmWQfx8r+cpmtPH658AGRIdyVySqnB42FJ
bcnErdCT4F8rehSfZcc00XH3wGsJjSiO/doWl8xH3suonYVGWd5aHoHU+lXq1IT2jIhDjAHZu0vc
sVEkPOnHGDRrguc3oQLxJsDOBEm4jhWpuYs3BMtwsfn+MgtuB+gJHU636ERHtzqdjYYQTqPs4VNz
bHxCNzvp91bvGy1NS/M2bqnDybA1CUFwbjNVYqLWwPxTVMc9Trv/vZCjt3NHFhwsdVFKPzLZ5lGM
hrfXnkn7fqDtWAtgzSeFUWi5Sc5PuqIcykf69BqxzBs0UaFnX6fgtdfJrF0Oeje04ABRYvVuG+eV
luGuBT5LqtABjXPyseXhig6uB+ZpfoO7dDO3onNJ8QfnStaYYECzgqMqJNJ/GtBGj0SPj4Y1riGI
VMg5V8rIH9fob4B9JN206j3tBQf/YzqnaTCCyOdu+/r6+gtvck0xr/JjfDoIu64YWkTn12sKL1F7
nIdYNtjQishQLq0ooq/zay8w8XAuH0uC85CmOX4yCidtl93aigGUJUHjIiSx9Rkx/i73gBtwEX7x
M6IhXe7fcggMG7dkBKd5ogpv6Y129xRf5jPxbIFfOqeC6VjXIG4TaG8Gu++R4lEXvFSVhAfrll9v
RIRhR56n34KRHdF/i53Vi1gbCauexMT6VbmnT2zLnFGm+WQTtBjOGXA7Wi/LQYuKST0Mxr5jf3qX
XUoE6dkecUYjeVQpRRgYLv7493NRnqv2UKEcRzmsledU61BNaLVg8PU75J6C168c4XNR2OK7k3TN
4NyGVb2+ENCKzD3sxmQ35ZvPj7nt02AYqtsx4NU35iec71ViVa6YXuy8GfC10+eOpdrQCDzPTZWb
VG4tPS1KI6Gbt6b1aR7X4A+Mkif6St0krnJRXHiIRA+UZ9ITo/b3pf1i2h3VnYbkiVLmmvLELJkN
lYfp+N0GvQirPKOGXDGZ0CbPciY6ZDPBSNN9+TLF86YlSb2hBhB43ANByV8ITun52l8vPz5vXqnA
PHZTgWY/BHvCgDdYVwumZRF7dPRImV1jhHb0qkWOZn0VvDNRivrmEv86qgZolLv/1plGvxJpOTbc
RW0NLDzNSvkTLY0J/vqPI9LFMVH44FX89V0ZS4xEUmTpx3qcFh3dgz/4FPSSETTFdpBgnwoMWOnF
Ptk7+qGRf+lpz3f2lWIxDj+r76YZMV0qlgrhiZI51+p09GPYs8aYcpp6gdbBe+gyZq5w2owZyvOm
VtWoOyD5cw87jgy1jQs1IpNIKDV5UCQ4IxQiy1jXhvbW9ET37hZJmYu/S/zMoCPSde0ZAzbvU2U+
DHowk6ZRGakj+8vV8F2l6lTa4aJuHZLdp8qIYstT4b1TV1aIzHNDwtiV1ZTMWIMBGX2z+npY0T7N
k5cQBiJUtPbamAD/sq8T8+hmLoCL22tRT+bmT+8LZN/hGW24Fvl6N402vljUHLmC6fAMb7xKd3BV
QVzvgw+oLP49Or2QwNP56FDMQjy5WwHlCxW+oRW2beSoGeT6LCZ40NRg0HCRDFNopMz0x+W5Z347
JiXd7PyjRjnd4AVkGa9UQUD6/pxXyf7rMs1WPuw2+V6RMPpeATINzkKhC36TAtLB9cx++3nHT09F
viWSHh1bQiGBGRTDbZltQ/bYtCh3YzbEdYRq4V2qNvxGrlqozswy1scFl3fUrqtUytiFlIY2Plb0
O+7+mUQzlIytnqzCvuvHD0zhdP0DZNCYYJKzF0YdIcu+IK7dE+ZNqmjszmUCEHj9qFntAgaSEpPZ
GH+O+M7VNnpg3InBaPaHDqvssFAzarrEi3/UEno0CjzLaCIQG3nmsZumOFcCO+GENt/MjcQwS0Gx
rr4rGojf8lTuVjUm+pCnWWiRgUKgDBlS5UGrJX+oGMxLWrPnAf1/UnY8Wf75S0BqfZIDOwwigE2j
dcrsbRotsNNFQAr9bfQMa1HigD0CydD4HDTlaD/BKw+T1hAeX2kQ4s6a0A/n+0CMk2DLU+654pnI
1ChM7uC459pgUASW0w0jgG9SzxkyrJeb8E+9ILdduZE5DylfUuCHkiaFicjJnu7CmsgULA2i3oaj
4SpvOckozfHxMCS7IP5k1HstUPDcGRpnjNxh/9hFdZbHObF0T/yLjpofyGyrNt/aLObVrX4cVkZQ
vH9w50Fpb5x2d99H+WHNmLxzQpsfr8lV3iCJ52x3WK/N9NzlC5XLLWAoA6K0FJSX73YHds/lceOX
t8mFWLJM+qO9FhUDs03CwHS7kOfo4v6PG4qnjxM3G96cOw+2ZtKtD8DJyLJY+PvXwBqhwVVxaj5w
qtm6nl6smfOreRnmzQp1UD0NfSom0ewPBQkc0ZFynN1OV09m0RKav3P80kQupwTOvgW2w3HO+hZh
eoqHoIuyQrhAg27wyVIpFE+viGqEUlxzTZ5wcoTfIrg5CIXvr8hxGNeeCmfYGHWtA1uZ0STu2LVh
VziVSZbEfgUvkUZBKOr0mjQPfybtpXOvOFSufyqIMDB9Z/1tKBP3XIz722pWUGyccnKKWWodTESD
M3kiiHx9ZWRKc/yLnGU8KSLbllF6+JzefCi6JkuIYFQoc3xPsvC1b1XXNl5UF8KkuTtKKAlBDPph
Vl4b1Aupy5gX8tJpWgsJbQYhPfT2mN9UxVqL6VvPloSmsHKSTy8t9inamPiRLhpXZiAtqnWCHNbg
Sh8IuOao9DbSpsRkWrOjKhYk3b+l66lFlQUoWVqRJBa8JBSYvX6jfcOh5JyXCjYLZAxS4i2XObTl
AcrNGj4IO6B2Bs9Z9O17khz7xkWXWo8GWwacjrXTdy2+Nd7fiAuwcgCgLOjEkWFwSbBudEI2hCA5
pXD9CXwqFvZjpn2M/XNVCX4nTmSt8bON0Ax8KHzLBpc1o1Sc8Je/QHtn3TPznBHJ5eosToDFZNRV
O/kZsC0QxXxrfrhQyQCwDOKD9w8Lvw7+tJD5siIemfF3MwO2rn0Pa1Zp1wG4xpqnl9YVq7y2rII9
LexfFW0dAo0ON0YhAkL4OElYu1m+dWX3K6lP1TqrtXIM+jb6TneU8+Dx6ib59Gc2O4zbVPZopnpr
C46W8h9AHknZw2Nd6NmfbKzUIkZ0E8vld6vhO4IQ2NwZ9XAmgaRppStqw/+CMb5gcoNfbkXzOI6p
w89+kWL6/Cro8887xRabypepexSnCZlc2a4VpENDp3M+lnvHrB3cdRFrOL4GE00awi43L/lW8k5n
ofYHK/Yj3psgrWL/CF1UEndib/EbiBRt8oTcLzGzREgt7xb3aqQoDYK+kKVVTT0LbVDeChs4PPKK
2t3vbKRp0HUXyErMHJs3w9i10Np0NtUVzFTao261lCdSiHJamaiY2c2WPDCr0V7D2ycAnLgb4AtJ
Hqm+fEW3ZR/fbJFrJuwI0sLG9D4op3+Bo72dzAsO86nLqpNlh7Dl3Xl0BuImcFXq/JKQ3kNO7ekj
SmAuxzVVDLqdHEl7/tCY3KH0O4uwpBqfvwNKPnfi2pQ5a6RaM5wt6TAPLNH/h0xD7N/EdtTrPfkA
04kPMmzmhgEj+pZIN1s4hutPDoFJNA1x8sh2kx1Ov3/26K0mr73ERuXUnxKeDVVAvfVPNnLZygJC
dxJoVbmBxb+426E+zi5Z1hSkULq1p06CnMCPbMbeuLaA1NsvoxNZXIuln6eq7PpwCB6caKu3jvDm
9w2aOPT5KMHD/bRqh3MLUFI9sq1O0WgBs5fYari1TCYg/rK8z0hFYpx6HfqiQWr7404S83eZLW4U
v/M9zVEswAJ/54s2IODVuD6ei8+OeLn53KxlGlGQ82CJVprn0y5rwxhGR+kkQaapItt60Y1SqDhE
wNEiOZe1H11uw0P4aRNrcNUPYK2+f0BOi50knriTJiv7JYHfp1aePkXmib0xjmxRrScU2aVNwn1L
sAhD9fpvc2m8PNxhumFeyeG+7l/0dEk7RqncBdN2W7AZWoQqHSMF47nc+5pXDX1wX/0iSQFkgQNn
bcINegxlch0l73Tjy+ujcwXK7ksn0p44klhS6lQtvopJq1/WAZbQHUCWlt75ML8qpY3g6C1gIMan
CaDhu6P/7ewrEX4B83M2FOAerRxVACcL5rtaR36qgh/G/1n0MqSTa9XmZrO7XQGSe7fGYr6oVjv1
rSVeb8vhWyLWFDvT7Ns42ttPdkrwuJN2nCH2h5kyZ4hkS1LiiA5OhNJoFQ6YtlNw4VltkysLmbaQ
3bPJshdTNdklNq9R0vZSTWewt4oJSO/sIIgcjaybhcyOjUHtfz20UyAI4MJYBKYyRfVn2nbvimCK
xxurPOnGXIcyUWwAgiPhsPT/scOsUz4/GgLW+xHW8LTcaQmJcgbnsX2fN/3AM1XFV1P6EaiZUVbC
4iItrsh8GxurFrxTHjRg43A/QIhsfS4azX66iEBpN41OblU/ixLKaDv8vsrzKaE7HmW33rOaMpz0
2NfCzRY9H6bB4dmnklvHpSFzbGIJtlvkZdiLYqTHnrUpYrqHldsBCtnu3IqofQJ40guRBLxrunpy
/amJ3B/IMaJaiQle5JW1VSCKvNd7L57iioPQ8MFzlhhf4y9WTMlLn7kGetOcttGmS5PzGyRy+Dp4
vi5iKaaDND0qmQsd+cF5eLfAL4d+6RnzLtQB4gGJPzTb6H+FYWAs3QCFUZrzj8c+sCGiZ8eiKPo5
5NrgdWAND+esZbrFiLEgCvIRHhD5a8X4G9xNQIqVcU8ZKZVNA5poQvdu4wnFFeCJ22hsqufhqu87
5PqeCMEVWSWl5rZRtXhd9MBlnWerO1Adr/rI5D9Tyv2UgQaOtZw8o1qiEl2eRieRqar1ysUNWA7t
ILqzPuNgaUtIFmviMJqNVNRFWEn4g6B6dLgEwoalbgZjU1gFFkulG0qYlRu6pHFbf2f2AwFVr2Kp
EDB6uoIFLQxkGyJgTrACk4H+meMMndF4cvDVYRfJZyERk/wfi6SiZ2PgL77VaH1Vw1rMJmYOXkvU
Ix6OcCA6bag4Tou71g2TKhIz8dBcvNtvIdCnaLvaCNtVjEStRzDoblpsH9YgfXLEx2vpBa0a9rdq
QWPPqS7TMO8y2WjECNe9JfF26xeP/6HpI1r4CGvvZBCTELDZtD39JVE68C5U733Ryd6IHhqXhTMH
SC1ArQYqQnpRyHF+R04GjSJVsI3QD04OIturKynRzWL5Mr01AthGu++QRNHda6KeWRFhDsoenig/
foSintsQP8oDwONaTjdJUcqYgpJeaMkruGuPyGpgVFF88gJr8NQH6WTsqfO5CZlBy9fcK29OW9Pa
V3J0KLr17ZKGn8SM+K7MQImJmuf7pDEzWBjWsmkFP+j/HgpAggjqFxR2IjRiQLzaB1qXVppxSGQB
2nxlLKTwEqBWwDc9etR83E4ZuguuTYQqbPLg0KRUu0CxBJzyygW4EmGzfZsSloMiI2FlkaHK9Ty2
QruXlas8pPCmtmTGntFh7vt0DiTg60p9K2lzYIbCtJxBvZ6rC9MB5MH6VEMiWuAY5SbFaf/jIVjK
Nb/rkI23ncxqGIw/nxER/zIe6uTQhg7PyoOCoo89M5MVdQr7+M/ByzGQztHb5z6cZHPDQYZZ8Q6H
sVMiz6WbujTjCKjIURsxzM/Ey2aLTHjbYx2xWEcYFO7sxcSzrqedCl1RNq1F4+VfiX1CFAZsgnQW
pQM7UmRuCBw/e5F+sGjVxSKl/xuw59oqlyZEWejO59Vrtw82BBKNww/6pHuqn7zNouoHG4j5GoxW
ztwLvAYtwNmfHQM0DTMEXjOCkBOE821cFsn4P1BYRe/hogAnhN8KAIUc0ax5IULmot8OotM4mYUf
/fIIPh1DSKl8j8j/d988k0/JNNzMSaWvZm3dmmexl3k2ORPpS1m72GaR80U/MLNlMHuaST1UtGgx
1M/TlwLyduAex3F1HGah9QxVuflP8Q6IT57oSCLwCWgXAot9QALzXYJ4IpMKG9csJn3eWldh838t
GSJRXP31kGRyioXJjUDUdIUnXDVwBRsIMg7VQzIVjXD+E2I5rju+iqGV3wEwrvlYwCZ4oLGZBYvl
1C4ntYHBl6UYk4WzKqqhhr45B/txJsRTlBp0B9vklZOvAiIJoqwbgJ9mZzFFGcm69AZySgPDcLzu
6TgM8w9FooZ0x/xCRIrd6cbkYVp6L5+icnolPsTz8tmuGUs8z9HjkkiIOUIQmSBSl69W+KvzXVXy
ZUhdLMsWBaV3rrjNpRKF3M/lKnF7ernEsXBTcTAJlCaa5a0c+2Bs8ru0eIsGji/tBCSXI8aZFbCR
LQgm6AmJGn2zSTyZubPkbtOuw2RqRAwr1kHt0NTaTdUGBZDSQRLs/cAccR2C10O352/krjiTrtiR
QBwcZsMT40+FKI+gPCv+dCzcUe2gUCAWE9WTLRQlTXltypBrSeiTi16u43bBejoWTRwRxKNvzOmo
vMsG0GSeuDsSdjl9halfAC+2c+tQR0/ZFWuX0wOZCnazev73Ao5L/iOx5uMFMx2z0e7EeOSkXV2c
+EjfFlFeJHV4vtvW98k+cvLjk4cidYOnnLz5YCoxdzbjm1IhpcWfTkeeVf0Kr3I1PmQ44Cc0q5sS
w4J41PtrIILDvMynjiauwj3rr4DI1ioC5KTyjCIh4Wa5RuAfci4A+FjXEHIFuCS6203iTlLE0oco
Ldc0lbIhz+4i7YeJ8LSpehtQ4baU0CLySU9cyqzxwgKDNRMLmlWG647O6djW7rfGlP5TBSWo/wsY
4Ukt+zK13hPJ3n0Ce7RsiJnc1A025cwHp8HwMnOfRLJaTQZlFy76oX/T/NgMdgyulDHnps0wFLXo
sQI21a3hNk4p0U7KFuD7JVe3HsoWddOuOa/SQuEw7hFsEqgbNdvTzACKLcn5eqW0jRLEziXCAHmI
nlFu5ek30uVzWnYZiYNkWt8UBY3b/O575f10rLUsqM+NsbkCPYd/kY6KFQ4qoIq75hMVqC+6flKO
YYldqlbob+toQDHgQhnNa0Z90G5Pprs9gKF+UUQOo+CpNy0rB7mhReJB3B3UW63RS4H6YWIP59F9
wXiuXxerTYpwwBpEx32zi1N1YU/zE/X6LAbSvoyLRDbMHUrGPn+OdBpN42WG8ipdbbEhTsSNrhDn
wthUx8bXMVK80p5msJHEEixJPo/AQRt6J3Lz9039i5UEgZsl9h5/YvCysvoU6835RFr8hkPQurzS
TdajRfzyLwh6d15sxXx9ZoaP2lVMWhnM4ACMkdF3uN9gB3zCoBz6OKQB/EHaUwJLQfTqx+RRE6R+
FzjWQuEprHANiqj2bTy3/1o02xAgs4mAlZjg+mNgMIlEHaT93s2po7tXtKqsmrHz3+V2rfpS2uEI
WtAbMqJsT4dY6yF2MqYpcUCW10MqGghoXVuE0muC2rZlSdRBjVJ0C/e6gzatKBVB/nVy4WkoZrsb
4wY9Ea/sY8Z3/t2eWkanJeAm66lv9Es6Gg3oFIjE8mbYE9p8UipwjrD8n4Jgq2a6cEmVBhjBMxGJ
88FnjoHcvjYwYqe9FdTn9/RdkpoBT5UcfrfrR2wacYNqVA6U7MbAkkiCvAdDLbR2rt8BIpN2N4mt
qPl55RlE7T678ur+agTLTl9IeIgrSY+lFgspSS7IMIw8piGxG7lJv1eHmgLT267dFgS/j690YwM4
L8cdMuiGzQF4sROXcF+ehWTqHqa+vzad+6HfKom6DTpPN9Hguaw8x1FJMpPN7tcKkuMTMKPoorNP
Ta+UBGEkevEI5CmpWONYFQrymmev3neByL89d8G51uuDSFHWeDcfju8jKV0w06gu1U9q3dMF79U7
bCg7L/GI4sdNWAcKkukoq7YskV/D9OsLJvLrIVbc4UEjdhUMKcJ0XetFBojxS+WF2SLLuSeekbft
fvO3j8DCsYJOC/IZ1snDUDUHbX1UCCvG98+TG4UWDtwNBkV4WD8he5GbWQ30kYEJ7OjCRFi/8qxD
X2v0PEdqna7kiZUv1he+al777QPK6OWA9MGtthUuXb2dcGBSuSSWrm3GrXn7pAcP80HF2bGoldEl
x4d4l/jKBS1iyELsr6Pi/bFczvrTqs7I8+VwVzMF1M/sFBhmCzOstWWOwnFbR+lFZc49SPZzScPe
2C/RmqjASgc45iMt55aGoWrR0vCIYWCWJPRg0fTC2JCHSaSfSwJGhoDKZVbJ8tvt6fFsNkhHR0tv
QZYmc7z8BpPOXGxq11MmGKSU5zOpNgByBILa6iJa/h+yFJIXCw0DO8Ul8miPdQ+e4bH869H4e81Y
ffwKs9dM+ifP7kB8Yd2yxuHhLDRqWUBUEKDGeJfZi64uRI4rvX5yv8y2zg6SDdsJ4BWDbQv3Zqva
rPNCSR97SztQbE4Tg20+06YTDafH6UdWd3iJc4TL6CmXy6ht1RqYc3Ez8FIJkykyLUv/h9X9zdsE
vHVh3B0fhfQLNSkXi+F+uw2RpZ3JrhnAw3zdWfmvWJoNQxjKvM26tgjsPyFfjnJpuUy0EpmQs31d
XAFljtyxod+v6XfHP0RbyNoZNuB15fjCh2J5cV5OEyYfGDX5U9d/xXCAq2F6Pi3qnFX+tScAws5h
fZJa6/YQmGTF26ZHSjNY3SF1WmmNuKEmpYtYykieNfi+7oAiHM3IlrNrqPZS0quBiFfca7GMqJSF
eM4DwwWUHmTPekW3BpX5v3q/D4x4QkWd38+5XTackFOw1v94apvFXfj/mDrtd/XYbFA7JmFp16Ml
4uDsv60ZcAXaFfjo4ZNdhZhK0TZ5EhYZe/muaM917sWKzNPVqtABfFUgAxzhb9a0SAIzI7Fs98Ki
eptzAMExNCQxNyXvbUe6vKuCpgdLw6q/tcpuHPYhJxxHeSLr3+IMnoTo/X2wXyNs8ShJGKQVwhX+
h2h3omX3RJXXXCHzueZkXbS18JX459AUOEqUxfEkhU3VWSZlMo+8TEF7TtA8Xx8ha9AoR2PhXnK/
EUZO+whDs3szxggP78J6t0UkSJrTnzq5w5CEMhFHxk954k00VPxONO3OqwQKgMaBeaylV7JGbP7z
aB3lD1bW1hPYDYYAtONNnU1+cH7E9uBMvvLqqAT9GgOoPdUazvVV2BbLLwTcWe7Bnr/ROKCGDTHK
kBJjsSWC/Wmy1uRs/hxFVKbu8ETUaswLTL10M7yZP2PKGIZ8Noz7uIcelVSZwgOnHpr2lu22rc1r
GnGeBy8oLnc2G4NCFP899C1mpilkn4MwbqXR+n6GA1qx+2PIsqjsQK27lR2HYgwHv4CKnOfubaZw
UxWKooFNz3Pz815HSMJGNweJrogobp/VVjrffjXDqS9L3KV12smFh5yIeFMaRf3PyRKoW9EX0kSJ
J9fXa2W5VzUrfNb/LpiK0+4VZJ0uQNzkqQLOmpitVKgbas5W74xEiTP5IXFdVUkQUANzpQltzMX+
2hbXELfzBW225H/V38C3uYK8+cX08cmX0Uyo0Rbx5zfQ4USViPH+OUF4z90xRrl1y/esDmNwhUvN
vNfpk6HgDB7ki3KVz4rwdlfvNwl1TdjIgzNLMSeVyDeRrbHUocPIllKTRVzGIoP37aUplhBt/Dw+
VAK76AecMhkYl9peJgfPV1/go7fOcK7I5GN1If3gc+Jok08IipwPjGI2FGLd0DZ6rhnqfTr1e4vj
tIXgehtMyGTXFuzaJ7IhIANTgJ5fzxUcplyoLcNlm0ZTnxqlrYpv86y7uqt6yocnHBwfuEij9ERj
zk2qI53NUY1B3faNcEyf8TGhVu/Y5e0Yr+EwI2hpYWUcDFsU2A0ynwWcK2OvycEoO4VGgqK4xT2Z
EGWVtrx/t9+ZrUssrRpahYO9z1ca3u+EFXm5aXlej9WUuFqkS2mnG1CqUZSbq/38yH3QszaK/mrN
3h3J6xbxh5gmyYeT4RpMK+lAuLR1Z5YHjiBMtXxTYHTN3PbCe+0P7O8KbTxmtru8CiHjmYGGQpgx
SIbi1DqAqG8Bg8SuPnIUKfQKL1FvV0Q0Jo47LNY+UghoZUmya7ZyiQtoTzzys01vMF4yvof3ex+K
Kt6oHEsO0RVxZhEHCn7f5Z09Xd7dIcomVXSCjfd5WUbEq19tuZkg0pcIvcoszQ/sjUD7kp32WAM6
lswCk7pdb+Z8P6G/zQY0/E68/NfsNBXN5dyVDFezKrLJOIaoLamWQst9XxjVtrZwLPkQRWhNogyT
vrmX8XUX3WkqKj8Z/bDUOIKdbTI8+gF3t+I+Wfn4VM6l1HpkVI3NZzkSHJLkwVv/dLEHlu173N5I
agPj7ZegNIMSEVAqnKRDmn6RUH6MIbhVZT2LXXapNYxooZ51Dp0wnWd/H9oWQC4ZMPvRBF1ZmClB
VkhmR7Oyt157crss095VnH/LXF44p/2JHMQRc4duf/SfVJrnDz35VH3VqySf7GXX9de3dXJcoj7t
4Oj9j0vBuvaXlUcQIXLT26eykxZ7viCp7a68jayxbLGSTymw1nVqmVQso1k8o/jVoK0RsSH6z4ni
QCpia0cArZN/Vnzn9Ky8HcjjZOZ42+bF4rLm7nHiKTI82mWlJjg2sHiPTi5Y/feGF3aWaAUEnYg1
X81R/uOCKHQsNwD8LpfqPbVqfNzssVIbhb7Vp8UUvbAqRTeieaI2O8oSx6btlBwiI2817o/HkqCC
0w00UIJZ2bvqcigCXTgk1eaZOd+cgJGFa483Z5U4pu6i1zH0DrVtG5cbG9FVNSL+NtXXY+8MEbxO
Se9a5tCv0oZRsu/hoSySMfFWIIrNdHxDLHr0fTUmDil5GVapX2/wPBmV+OMSACCFRYOgmcl1oxyG
Wkb9LCDbfo3JpqCPJnwUWItpR1RzQ0yqTJlVJ6m8CQWzdonIyjPtQaqDo5yT9eYsV0TwkoatGeHm
oe68Y43KqSi5rO2eg3ZLSi4G41oDps09+x9CiUnwqZISueQprSmhPRsKxk2QD5LQzSL+DY9xq9GN
z9/Q600xGENPJrcQgyW59aNqevbgT3f8qJNwVE5B/9lkFnqU2fZFvdxunBSCLDUc8XO7/82QuFmR
RP9x2qTeeZv++NkwYuzEwpu3WINze/KivoQM5FIA+5spycpX3uvhRrcSReSExBB0ygCwATFliYnT
8GLBAoaqi3KlgjdByTmi/+SZcEgvqWmOPpDbjlnpcQoUUsJ2AB8TmP+uWAUGEMARHwnfYiuTrgpS
wzpjMujGggUI1ugPF5x+Q5gJOMQmUgSpUb3dJTBWthWc4v+x2qruogkbP0RALz1BJRkl/mhKDV0C
45pdX/aAoD/heemCwjPsPVGOvW0N041TjHgOdeAb98p99VTIcdEA3JhVnP3pMjAfPE9TYvdOytnr
pqTK/9mnrF/74j/01VJffAvJgUbmeuyClZbMZjcsaCEEFwuXp+NCcOP5/wvFgvG/xcDGzmHGxiXL
GE8XZhMZDIjZuAs8QvNrkLRxfCWD8Yu3Lo1wdUi3sVdZQnQmCuE9hgcOTnZivOEtYtZ72DDwM5+0
iVG/69UqZql9BECC3sgjpnlwlPs3pLrONCRJO+/i0YdEony+jIQp1dZw7f2eYLQT66LETtz0a10/
MfbaU3jsgsQEbIlBNsiVdDjhNzn760/Eo9lIneSgsrkgebTbk6/MUkX3FPYgkLyCowlPexq86d4k
/Ce64vYCgjvArsc2p/Dr5BQJVVH9GXjsOoHL1VaHszFB10gaZazYkYB12LGoR75j1yR7zvGCDl8r
8s39AtcWESmAKWYiNoEoZcCTEzzphmkk962yARlisjZf/l0DMxhAmXs3wchh4lxL3+bErXYe4Rlh
/GjK/1Ro9TM2rWB48w3mK/QDxoy765HqmoofSd18DyXL+hLFzJM0W82AVDWWuz+5ZWOfq9d+d7il
0hX6fbNQI6Nkn13GFm73rd/8WuTLRxdzy17C2vpX3Lir4fbxb+XIvoLAC/44tGkrLfSukbzHmyjw
uVO0DBr/rholq7o79bgnSZ8ET4vJBUyvebV5Wqx+JjCTVD8xyrhlhLqC+xDwhkaGtml7x9VRaHqJ
k6nHgYPENQ9xQkZSUbGv7FqlxayqdnImAZq+ZPG8sTg6zr44WYCZVTCVJu+K13Ej2kEHsavmXfO5
pVpMERucKtQ87tmuJiT8SuQMZ3oUQ012uzpI5MDVd4ZLVcnTH0Ou6d5Zfc0jMBcqagTCyb04yF1U
Q2LyiWFebLYuQ07AZDIxWpDXS1nqcSkvot/Y69AelroWNHBzRH7UyS/SvYmnSc1RVuvgp6V9jHTu
cjr3JQSZuOnEmzip9II9Ab3eYUwGExiwkqV3GBUJdqk1jszlm0dhQa5Nto5+ebwIRItGwHs15aPS
03KOS1uoYlHUPaYEIAKY4zqViOyCbBBbiqeMvm1Hyt7bpNdHB5KALaXRf0a0bMYqz1oeyOgg/0ca
QSZRrwS1LS3DznVWeJDheuzq4zKpcsBrRQwh2/7ldOtjG2O5jz2WjwucGf++27xkK50ziAIPGtQS
wcwQkcFdfU5es3i+kb5Pz4PkOmNKh5XXJ1knV9lkgR4clKGqoHTcrWjydHmFOXyCjdeev2DOzNwg
6KuKYgENXLL4tQY1g58FDMt7mHYoUUScaTZUjctYYCsZ2DKv0yg5xWBjsO6nvB8Hc7pwvlzbjXM/
ynwwCqgseSs9OWGJhU26VQslswiDEN0++bW+PejoT/hewFM0qZ14Vs5Z2sDNw7faJZ58auNgxQuh
9wmeheWUvTNOkG318IxeCTa3S2TZ5wGm6lgswBNC9pWpORDT4DOTVxv7EC/hwuQUiO3tVRujZwcZ
9kbSt8G8zodqnoscwpAuOZWmNB0TP0Ae9+rvsX7DiFiBJO/Fhd8XCS4ea3KORhoqeSsY2E+15GOR
POaa6TDbHRZVxrM1MTn95uHai3s+TlsXPtFnnWnrELBiIRdZmewDV7cfJLtazF4waVt1WPHnXss2
ucYqIDtIshs+E3Lw8pjZ9klGN1bArCp2V9sK2rwVykkTwP3aQTJj1yfm9WBZAMMh0KeQGJZ7eZ7P
LIi4ocI5N2tZ5yjApkhyFq+O0AqWJda2trCsVvJ1b1UmAw6YtpP+syh64ENIiUs+ZCo66ugY49Ow
86X53x77z5552mNckedRHwLCCjSXoLpCoKcnetEYrlTB3U2Jgl9EcE0892fLTb4HD0IrpSZqP4UH
LxY03P44zQy6Vm62dAOL/c2WAhkM/XPzQ39NboQK8T6viQweBXAEg5CuoUq0ACuAFybsfjgUBtaX
+WzoGvPJeQeIu/dmxMZueJY6wOHgUd76hK52swgY5sacui0tHD7MfPM0EiOEdXMQ8xp3a/0Nu8yW
r4PZ0gbiAP8nX5z4bV3LE+1adCrLEsx50nHtXTF1E3ef+YLCIteqoFQr3/8/+3KxKr1bazqwbT39
czm1PqUQDyXIeQnoq+3lPo5sD9dwpBBsHiepYYdJTAQuNy0CF8Zx18rsNMbUBzO3W5xZV6efn3x0
MPzyiwfnFIWbo4FgH0YyEfTU9jQe+icdjRLYX3mPIH6hJqwoyDrsEAznKO1L28bHU1EwftuXNulX
hhGQBj+y/9EMVNhO4rX/xFxKR0uvm/0Xah9wbwtBstWMV3hHBmq5P6m1p1sEOJOdX/wd8CsbGDDk
uLcEnVrYqpICTLrSHeq2COKRYA97CBc6c0eADUAlzKIwR6KX4PlQdg0TLqfr/4iNrhnDDCpCXuyT
tlLKu7rwQ02fF21F21n0X4kpovVtCxvY5MF31iUia7COkUM4iEJ8qCz1an+MbNjbwGDKIOHDbNa3
T8cOoyB4ZY/GOVP7qSTOlOrISgGRVKYKvD/wYEAaiiwhk4+I7Nn52a7CbPANlEdn5gR7pRJ7H+Yn
IfEB8+Wc5zQDg+pjSVEeoQ+7ArDqErkiXY7usxDsddCLJi+xbSiMJNc8RblmBWOuKwRMcGEkkTHj
0G4+LEFIbYvtZKD2cEz9pNrF4Nc4TATOpOj04rNJxdZW62J+iUl7N+9o28L3344iwXPyosaU/LwS
7Q+NkQMMkvI9NM27m/USezHnD5LzktcUmX+Ibr4yi8T4fOJMBwIyrZ8jS+Z/6hZBG8/kx9lIwcIT
5sux26kvDwzBHGvGG2pojtFszPPA0FHF8IV5Z/+qPNEjHTExAwCF+BxqabDKC4f2qYKWVf1hnzLT
7M9dytPlJOMMx0R1T2baaPpVTxsfG2RmLZKV19SgMlDF0SDbzfAwYuMKiHWQKP3plCb6pINisv+D
vLH8x7TlRYONDJw3CndW5WY+fjbKstnlSICUynj2q1nt2sHUZ+ddigYhdtY8vPJXu7gs4K+cHPvn
Gvry7uuWRbWFvDRFHnV9R6QZabCHSnergYHOIjHSnuGkXA1SCZpLCCu/caqUjXaF7SUxi0OXbRjI
8iU6npsDbI/MZFWe0yehtZzlpTyWDLFbw02cQvylRIjeUIEuMUvl9HZETu/BN/DMb9j1dcjw4Ocs
KRelkn3rCjv9B8kuvC4rq/u+bJNG8o5JB3XsOCcGVV3YjcN1LOe0D5ICK6i/GO8OZNylygBSXcn/
XF9UrIBllVM+VT4m1umGN8j0WWxrGTQ8H2xWl37Z1CpCMylbNZw49cShgYE3W4285eQgRcSKUXIS
htruRbMG1LQXBmRvqgqswqSfxBVTBHs499IBgADhurwmikdMxFeauv3PSHGFj9X8G/7MFPO0xPpe
KAmTqRCH6LzuFCMCVlV17XzX29RHz/T4XBGOUSqTqb9v318U51ZslEQLc6WsmeenB9JJ6+HbB2YP
KysqPIJcQi7Irb4OckMRcFzdwcOiPYqFmAH66TI3LFMtG/r8TphpKHDuUTM5EvW0LbHJQSQBAOKr
PfCyinj2RjEHIyyrFY8zGsYAM6lP6nXAQX7yEnG32bD1zvhfmdtqFhcI0EpYEDril6/g9aXkdILw
XmsjDkqOIVYeq28q3QTXjsYXNOoyMda66HB/9YXfPocwgvXVA/FMx/B6+7gr25XyPQ7OP2yKYJ0c
RVDg8Ls2jNDhEVemWegfAyGSZlNqZd5FqO4kmQHiWCnjWtdz/q+N0+jL7/6jNfQiVwM6DMIF8epo
OLVbf+23rkrfe0UdLM3GR+19Wk11hauJ+Pc/hkaZ7tRYXOJBBYcCj0qPt6WfWtpWGSgVRjUomqWX
9TRR28i6dz/Gf6gVfqn0eMA993GhCyZxllUjNU4Njk2KvC+mzJpU1dXf+PClrqg9Nay522YE5Doy
HD+toimSM3+DI4bWHgRqyi5BcZWbSRABUTpa4ML1YkcjZWO7IRDzbdU/Jdg/3Wqv9blIG4JSuRsV
6RaNfojfySP1tTuU6RGo01X7Y5ItrJsPY2be4UOypeTGHPTo6Yc3VbAUpmqOp9Yb4311JozxR8Bx
ixjLTqMoDT1Usk/DYDk1JA5g7Z7bgN0XMi8o44yba53DHqdIpa7JmYGwCeBF9NqmJ/jrSIwTa2vW
rKEJlgliv3cmPRb1Vv3uP0hv08TZdxSEO5VIDzCJVcR7Ukb7w9wsyaSKqWqjloGhW0ZWDjMGz3Et
cvx1eZ3r1vdD7FEI9B+TymheEXq90L2PL+OGzRrWqBQobKA7bmuib8yH3QfA738imrNHKmmjvL5Q
3gvaP8kMf8NF1JeEndVuVRmFChcuskjUIAU5g1tfJfqXc88PGZPlvBj7lzyjRwKA+YnxXgI1TN9Y
G+TN+oRjWZi9S4jxquzYeaq0X9+olZTm0Evvl9w53fVbB5YDpQA5L8rWOzmWXci0PM/JiuVJlHxR
BeNtz3u71Yuc/oO6Wl3njvqSLavnmYe2zMbheGNcxpsScKXPBSbvfbhAf8+Qc+X713w2+VLT7aIb
3TORWTVQgMFUWHQ9ZB+rz9qQSuO9fFsGRfQ6iWsaDTcr25SpYtr4Vf1Y487yTz3+x3U0uXBkUJsO
KCxO+XZkuFospuAnnL+pxUmIm+TLfym/YH5ea7oy+hjmndBsGJdzlOWorYqVjYToBxn2DXZSmy3e
QCQBg8fkBwJODcFaHRZET7AvUZ0/WRxainuDljXuItTu+b/qPBU1aB+TO14EdwhcCbnDXDyyKyvL
Efm9wwwQIO6iEhXEnm6TuFdjZwY5Jcjwqe0MhSIqcTLdt+r1hRZzbEsNXzWWdKauw1MDrJPFQni5
d4nGM5jtmmheM2b+aARA2oRSk3H/ih0jYGw0LdY5Mu7YJOzyrRxuYPKa/f6jBIdpKqNa1K5RZuDn
66CkfKPZkxgREjqwu9DGCYfnzT2Nyxdpv8g++gSRTOmDn9gf6Nwgkv52zvoJbMjw4L6ACc4DAMC8
F/9amPw53R+rQSLAyVuG8bmKhn4BdI4IOLP8VWq2jr3lfPyOr5ataud2KVrOaaYIGa/+Azk+qm9R
kO9vjvWKUxC7StJuvRQ9R1NwB3Olb7y2MAz+5IS1rjt2+5265SIO/IbvfyRk9wgJpA8nA4SX4/2l
v1tvHWBMRju3huE7XyoqU9XArG4ARaX/+2ZLC3ezXE/mQUFBCAvHX5v812q+0HUZBT+sF8XLPmUU
DMMJTJJc1VgFX08lffBu/7XcytHllA86St4wIsn3kGO51k/Gk3y+9Sza0Hs9lCM/T1ZRkOsEGYBy
C+QzA4DqpvVjk4JQNUhV9Vwr8GOPQ4ll2fvFblfnlFAcU+kRMzo+uKfXN68+f5MsYqvgqNGq1hM8
qfidFAow7SSn0InOiINzuxVrCxp4ks/S96LcKajmixNqYM9NwcQnTff7O0cem/5dLfxi0qJXgzoV
AW+NBXn0K6qBShuRol7U7RELv19WDADT+FQJypNp2LCifq63dquy4CrERgU6XuIKf0G3lQHDNe1u
BOGeF4/CL1hcHf7OgQ48DyeKt7TBkevqnVo3a4xJeUmaHZGNPkl7LIikwbppVI+dt8SoxH9zimhM
UpLiJ/BitGFlr8adFeNaIVyFv46qoqNWnvY7w0sFVseVaUEDV9ZNWI6TdJmraGbXJatWM7Goj9UM
WNtLdtBTGJoSiI4qxyVk7rby5YbRjhhgeUFBoIPwZOyGA59tlGX1n0E/cDA/60PK+K674PIKrLZp
Evm18km0pK9VvXaxw9+02jcfKHqYZ99clIrPWIb1kTy/gu9DYeCxzxsBLTmLYPF/EHrfKpUmsbus
YNLM9htVCZRRlUMtI4ysgZ3CXpNo40P1cAaB6k0yZitT7gBb83fdFGfeGG2Fb8HXxnBOaiiD0Y0h
I3AXHOnFOqYaGQ/xiO9ASS34m0IbgG+bFHZLXZQtrzriKlE0KZuc4l/UGObqUnVUirA7jLJjIspG
roDCdtf0sdPKrBbs1HMUIEvYIcMhKLdFDwhwuRBwxYMGa5Anup3WdbtKJjWtbSedXBBaE8JFYsWb
8p2xipbQgQYEytZOLLGyigCkczQNJW8P+f5xWKY+YqA8n9847waMOmP6/BfvlhM5sJh62P/iTAFL
2J+MNdF5YDzdkgrZ5cnzzyEnPtOM0cGmbtuxOZ4vKMTdxeb62dmBo8uBt7acLY+2PgOQYozeMzGZ
Uk6Fw0Dac9QknSfsYpFbceAnqUjV336UEiu+k0ppocQsfl8aNoktBEdbaTP1Tfp3cagv7vKz99S6
81fmUbG8vf1/u/K35MZXybJR0gaDbg90ZEoclBooE47W1yG+tvRhhLjcYFG/WqDtMlOp3YNZjP2j
IC51cgpG3b/r/siWSoOEbSrKZUrDgQ9yiCeAEgohZFrugDwE8VfogCXd0Ku0uwGZV9nURVBVXlIH
Rusy/HtyubgqrIjLpq2VWTiv6ouPsuuBbNO+QeyEIvjL7dG2irSrEDxwMWp4h8JJpuxH7g+rkHH0
9gPoCF1dlW5HIXp//a/r1SCV1i9hSyxLv+RujRFaMHCsYRNoLcqAlVVEK9iFwz7pafZ7xw4Nja66
XAZFGNo4XbdqGC/5yF88tSE1qhRdiOQFS+Bi+zeDOEvZ6xFrtqudocsbpRXculTL+FibTdpnBh+v
ulvNrx/v05+lVGgudNbrVTM7JcZqukxuzPsxFanxTc/fFq7AvNqsJyhmlnWXHaiteT6OJQNKEmn9
2UxOs4OjMzepu/ll72SOk+Sy0rnNlew7hXLVihlrStKftTVeJ4B7czaNw+wYIKvtVJ0BwQUWWabS
PDndiIKXG0I5jg+wNMAd2e6FMllck6EP6YrSS2tVtRbbmMX/a14hjlKOW8PVWZD8YtDE6qHf7YS3
y3iqZTqblR2Fofi6C8fpOpGURpTkbQf+oBx59fWjS/vCJcqospWe98pEJqI2QAssyMMlJmtPbKfI
mEkfzUFr2B2cG1c0gsZEzRlmAa680gufod4OdmT9/9rVHp463syxlcrjbB/K+3cl2Nnrx5Xav15f
m83GIxTUTDyjIriy5EXMFhgahc4NxKuTVJPuWWgjlaAfoD1TPNzHqorkwlkIK7Iw8LvX8OlMSCEi
bjln0bbYknwPYMVYTGu6gMlaf3PaOSQN7DmMwGwHBBuyh1PU/iVxH7b9vyqJKcv3j+KEbbkynTau
qvRIV3Y2l2Y/kVD7vJrg+C1oRNi6/OLP8cl3H6dvb0K1cYQ82ZQ9MNmw9wfx2Q9H8Ap5FPoZQiD9
Q8kOTWG0rl0tfVKK3lmGklREI5SUmVaq+FmIP1JuP4ed3qpJIAKLHJtEE4+QCiqWlk+b9mUuPCb1
jMUrl7hDPUu8xTOg8IcUYvGTiPS9njUMGFiRVEMt0zJgaSO8sg+c7WGzqfBADJhTT6EzbC2sZkXO
I0s1Gv7gBYuSZ9No8yf8DYpC45FFv8vzd6N5jEYE2srYuSIRc35xcbanbOHev6ZP3mB0pl/+7T3w
bbAkrOkhJugRNpk2nvIOyq3ima72oXlTxTl5T86lWsdAnpHFc01HJvcLqk4uLKpg/SRBQjfErtFT
Bv6+AYHMb/oxOyPt1tKYC6znxt3Ks8As0DEDoUH5HI/bzsqg2ZoLN+p1Q1qmPbJDPLlz1gYF9gBc
BStojSn5P6xkfoV4ftuU0m/+P+PDL54yFzGQ0U0TAsz9soHXnm80LeLG7swiJLZGJq8lK26Q8raH
sqi009kuwHaT02mMfxPmlV5IQBm/ixyhmopjHViotlWeEyUbeUrQnnqzwdMgMUlmOZipIy0//Fri
CyR37zepX+j04iypkSz01ynETxXcGyATF3fMAmtLT/HFIqm2PxDeDPTqzTbJx6EulB73bd5ymBvv
nkdheBo4FN57x1mgZM+CisGK0dsIktgNQzKYvStQLj2OQWdmSUbZq9CNxarwNIFNxnAQk1dzz6/X
dqZxaEwsxVz8FecZ+ss+BTREaEu6pOxTTvRi0LFgPvcGMS6uAUeORr3TMKw6rS6j/9Wd1lhAS8qg
AGGyeYUn52gZ5IHEcaD8HPZ7em4s9cI7G4SvKsa06S2FJUmVmIUp2T4io4z5is7D9mZjFf7rE9ZM
qbKDjSeeTj7pyyuKdvY2+Bj+sySAhSmidDfC5jZafDk7D1nt64JZdNTpFkuNn/n1IHSyS9gmw2Ra
QAWprWhA2CC+k4l9z8aXuSuQWatLBN7YZmBIdn62xrYLOXXese44LKYYPg1w2C2697dbejc4Ro24
w6+I0MKbPKNl+trhrNqqn54R2aweo6WPzlR5g7wk4DC0aULL4NQQzrKxksDGxHjWxkI6+FrNID+p
6FVKqwUb02p/tSZwL8FwzWUttHwIpaQ0kfvyeak4T4bgEZn8DVawcZG0+KmUzE7atX5a45tgYSDe
tXtXOKQJK6sBjiuAQ5nIvs+ebKw8Z+EKom/48lkFQ7qmQYsvYKMyvU2WC6w5gOzB9j4gp/2/k6n5
K2wvYiBmjCadf8NRyz5UWBH09xwRChArJhrwI4E85nMs0LD+rixb54NieKO4NGevUDyoxCvA3m8E
7yu4atQhYQ4M6ww7Y17yEcmZ40RohAY3iyFceDKtRInp7/g6LC2dDB/PRQtp5sbWR+0i+rCnxJhW
y3gItDHjkq/PKm6O9MynVti8ZurB4Ux7kQn74/PosqSes2M9f4RzaxSTbCMLIj+wBMb1QGLZqLAu
jdFilqlBISG30vw9eTQewgc8PxR+IuDR1xq0sP7kb8834aXWx8qQwKwpeM2/dcyJ6zA4j2+yluAH
ayMiDyfKg+qAkVH/yyNhg0xGbU3lHjAQGQvDcuTPGoJFn9t8tqampx24lrgVGJXEKiDpFBu/V4Z0
6f13X8SDiix/D649k9l8Yn0uo5tuuBALGvtWUT6cf6p80R77zykS26nESgYM0WS45ombE+Nv+P9P
8vHSsteBo4MTmAw8d7Bm64J95kVcgMie9y1fxDlYwDQBW/ZeQkreX42BieW+iKwPyTMKK51J1zrl
0mOsEI+RyUTMCiBzdbMiAN7NOAcxFajNbiPIDD1jqrKaZrgnkJPO20oej5px7ywArqijhzST5XLp
g4GHkKZxpsGJusEc5jiXtPUIaWLFhnGKCn65v3Q2GSEnCP/8Y043hLhRZLGr1z01LgoICk00CxUt
MS+A60C9Yp/keaBgpf10JArkw07mMZRFa0p/qJ49kGgxQrGMTvJngIHYcY1HgTrKcz4iznQ/BimX
PVCkAxxlK1YlW9JdjEHaxLDBG3sRKFyZy3U9f7JsG9BA6efvOovSK/YvKEqQTl7KYlo9fGRDQyea
9DptjsMgD9yLMgis1OY1IoqiOPzaB1nSdjF99sHik+Dm5GRyMPYyA8HrzYT4iR1Leuc3oVoWk1i1
bu68uR/0j4/O0itAeBzqVgXQFVQjlPv59IGMt5rZ7Z08+N1lHQZhBiCZk/h2JvoXNJ32KSiHq6MX
CCJ86bC6bYk2CJGOftKb3rsCLFnMphU2wbIzwS+WMKUJeWuxcRGGTr46OawHKt78DNKj+qrH+2xb
TO5YWtjrRYjQKbuOzQi/Ic5VHWk4PYJfn4lZuiBu2G3NQhTK0Y9Y18c8oWq9A/ms/HqV5Ug860cL
iCuimp1agTqImnFOjc+f9LkmQlvZljSWjJ577KIg1rXS8Ek98RaTyV8uAOLAGijdiUU0gp20EfQC
NYHkHOzrRvKXiROLVxNJAeYqv8s/lFygTwECZyDoap8aADYiDu6mgCkv2l6DzG4hYybBmnzYZeC4
fvQLPr2dioGlr9P4hz9/1l7o/ia2LkX7QTKIt4xTc2Cl+fMWUvRRrZDIZldecpRvWMoRPo6gfXSQ
yt1UJ75X1kmpUEJb0UYOPBBAIAff+YzjUjDbDNO2J5/o25mV9DlAiLYd69bn7LDQl8dmEwS7J+8X
0nFFgIMUIuy9fdkEA+8/kCOumznQpHndvTrxXuwLaxh9HGx527XPCWjfXf0mFnSBKCljqun9OQX8
rjSDiE39WXWlGOP7a0Ujo+5LpXicoL+dqAU6Z6RlvUaFGYkiXDb2csd7AiVxDAH9O7+xDrAcgkNV
VOci7nf6xR1Ui/YVAZPZP1+8+FqAvypiGux2l4pbKt704kZ+HxKXoxwG7q999tbgNNUI9U9KeMPU
BCS99U/bb9LTBSOOEMtjEYtRez/pNPmG9pCQuBXbef3Sl23GM8RT5o02jdASE1aj/B0/1AzXYpOn
CWI8Vpr3JtgkGOv+evC4AJjdC+SMw5qOflH31KMyWhLpkZ8UYMLLOEbVZqOAgl0r0k+AU9zflPum
YMTMGQ3/HGwVESWUwxVpUW0X4nuIJ8LQnJsnE8a938rsI1rOB/2x0OIREJPIrT3kEIThSBRQI4sc
Rvw0WiRdn2GyXPKVjsMvCukyFzIZm2JGVtslHLUtbxBcAvlpdikm4/aHl5gBxPRoJM0MzLee9Z/H
Ipi2Hg6vuK6PXkQVxpA72c+jqwI+OcpJx2lThO4TOf2gMYWi1GTFDtrvrEWrQZnYiOytda1nl79o
HP5vC85ZMe23MFqx5DT7GuZwFFgGkn7A8GCeDPkSsJhZQGMeSZRyTIQg7lhLcAzzVmSlwt4UjGvU
rLJocEPhBw6hxt8LXifabl1s7TBNpmwnDt0cuNn3/m8Qf86fn3aQQuRgWk6atzh3YN9OL3xcQWzW
6nQv7r9avDJXhfDWFj7uEuVcEaN7y7nHPoYsfBsaRGXgKFDmGKr9VzIqw7R/aW443r0il/P/5LdG
VCnU/sR6gy424ZdTBq+qeyBlSmsbBbGt+XMjd1apEAWUrCD/U21kJnjDQY4jvqoCKw/jTwqZbO9v
1/uXVHVBRMTGWvQiquIoNSkTJ+PVW5qtkhtRroc4bDL2K9dk3qikyLeen5xBI/5Yq0q4p1G/aE3Y
NLQzWLtpyBe1zGbQmAQdjetfrP1mjD1lnYBeEGupyZ893LJrDS1C61KoUBscrBYtldpJw7jbmmDV
1ZUKNFUn0d/mhXJfgFpl+cfCpPqysI7CU8dBo5QYzn7sh6wsrtn4YO/GUIOMMa804aeUrn50LD/W
04UA4FhF10G5Zkai7pPvFaKPs/HQjmXv3P5aL0FFezbEq8vzzYOpkBpnMd9HpfeEGWj3Mwnt1Z9e
edyhsMtilhbSgINxp5ylXrk7n8wF/1CSUJqso/Ndd3ztd3X+mjEv+MhXz96yzXfXS14OoMkmDqRh
mZNVaOAdQm9jO/2I7HSmLXNxBYamVcWASW0dU7oAdSqc4yMZ7zS2Z+WPZHJm4GwYr9MpNv54u7mS
QVhwgExqyo3KydO2a33dk6mBC9tjyE67Tpr9a12uYgHY68SqBL2Env79wmZb3EqAyeysa6bRH7fu
lTPqWnKKaR5obon7xAp8yVft3kYDR/PBi/lhtuvevycdJKhMOO5VIuhq/PMGMZvMfJfVMQP62dfo
/XSbRni2uv1efCf750QWjB2pKctKsZEZXvgsxtuNC4TVHvYxHCN8puDeRPXUAJYvV1KMaCMEEK8+
3RA+Mf0SNXVi3sCmcE8mmWjEDj/QF8/RjHqoe4eTKat1NmL7YVAY8gFducBtTt1VUyuh9a/Y/DeT
9btyexbAWwl+/FB0OlUP08sdmnzFojTYgAAtkia75/dU21hJr/VRN8Pub+dd0WoRzdqbK95pVCZ7
OjjtJAKxX1Fdv7CKzmq9xvQ8ivN8OoSPd9npLDx/NnkWq3yrZwj2sPOvjbZ/TAtXpwps7XiMukXX
osuZ9oGJhaqcqBl9gIZ6fSuwdKjNxfIxM0qVtxZkFKnqj0luE5GOJt+2JPffzCbJ+fXyKltj2exD
AHrEgA8L9J3bPFKG94Ecm42A6XeqF6dEcMBN7zaxd8NpQqGlgKC0eJ/T65VEbClGndLrSZX+LN68
Q4VTFG43ITx5d5e50i8sJy3l5trh+PDAgOFFDFSA9k5xm3d6viPsJ4mePltZSXZin191SnsWKOqt
jUOypuEA1GWACNnTbzI/4vBAN8dBwXqD1G2yBKOGLq4a9uheqbhmJwHnZ5FwViG0g23vx5XWGbYE
qnMmndnuEIXXWRxN4Mv3hHOh6EFvXH+XbzWj2nG/bP0/OnlSX5h+Ud1Ikb5nma6GYM8N5HTADun+
epktmbBHfJhtF3vvPNc5kiqonQcxqwr87J2NV07o/TAlrJtwfmXJNVw8Y9Qz8KTcreFLbu9P2oui
xfywF3/IPM+X9mFKG6XKbsgUIte6fRRt4z57YVuRqno+9MxSQqQwzHF4KAbPwEGT1BiEx8o4EDkZ
QIVPPUC2GuooCMctx7vklIhlaJ9s/55SP6i5we45vETOGNo6ha5jtN53FNx7+JTFvnr5NqghysRr
PhfpgFkP0LK7u+yMxmz6KvQ2yGS6UBGxrGpgpBBuTab6p1Ggg2AownMaluuJLabZPDVasV+GXRQF
ApSGZDk2Xmoq6k7smoEBX2CZrmaGmJXm04e2+iYvvfNknpwNc+FYy0Yn3Mp/Z2EanBUX4KSuSBEC
1HMr7pF/cDzmG/0uhQK3P8Ow3+DdorgA61gr5AfTaQkzyY/tLwF4dw5QY4HYW8EMrVlY4ITdFO1M
GiXuwTirJkHFxEoDVHp9vUsebBNoax2E8YmTjy8dsH39uENk4+16hPx0egCHYV4omxAaFx3QvGlJ
IjrM2VeZ7GvH0xpT8Z5s1EX9/pzyhR2RlsEI+XURrEgg4dyY065P71pze4NiduYpMcwb5e3k5+Dq
okTBoORGEae00XH60OJbTykc+6+fp38mSd733AOv1QXZ/zdeLsQHKSLXuyd3K6qnANp8rcT1w/cV
UYNYhGFXfmdc4KK1GcO7uJnds2IqADO7E6aQGYn6J100/03NpttkN5ytKcqX+cjVqTLvcnCw+hIn
BECn62/8OCNeLUKFZbDC4IdynjAPs2Sq5unhrAl9DpmL1Rq4FS64eJJ0X8jbhfdh6AQXJjpR4fMW
ZzcxvJx2LwEXiolrHS8vpNJRcehrC8VwqYUVzW1Fqt+cZCCsgv0L7BT3rbwBgavsws6BhIF3P7Cb
tcHLg1T5Cevfx/c9fp+CjBuHaFt4h2TaMqI9Sc41KDrg/B+geXjDUr57Nuoh5Rq3fFkc78bST2Rd
QshG3DVZ4bwsKk7PTC4mgkXGeA775bRPOnOhkX6p1MUI4GLzLi4ZQqF1V/pnLJ2CKunGyvkvcx6D
UVXJ6TBigSLbG67gTAD0uGyotCqEhQz/4yZQsGlvJqMbytzbmRVjHsPJXoa4nGzQsi1D5qMrYujl
GYnsQtoPbfRyIVXkWPrapSgzr13RlwDGUJYpEPkct5PY3oWiJfxMhCGn43CCa9k7BmnGKnaJvjML
NogVZgwkDEU1RWa6BjnUS7opCT7ZKsJ4KiqSNLJEJQSnm/bI2iWL1EhLCLh+QOtgBxZxNxOBfdpu
pyFvS2sAnAKsDc7HIWT3JlkB+2KgNr/enjL01xNmgJSsqwHrf1hQz9cPPnEeP+WqxM7i8quagQl3
p7bGhvll5ipQX1sxIBrP/cfTkFLSuuM4PuCz/KuZAWwVmOVsCCxlsakaE/LQePFsaweXSg3FM469
c4IHXLacPsR67CpOwMbIy9Y7LcYRvta/Xd+SQZIurIhAnhef+/wCHU0iblCbnAjfyANiHds84fhe
ftFdBQ5AaTy0yNEF5n1u5/7jTPEZWNQohsrWmTEPHFkuCN1535ECWtnStWABvn0IRmGomiSSa4ju
qN4ZOSGT8+jeaoTafB95pzcoAEb83EytVMGruPFz9gJpO0xGJoUPiazSlVD+riZBwGDXKovfVLDG
Z1hDt/l+WMSnwbdXuFWK/u/4H8EAFP3lA/pJ2h2XyBY1/WR1b9lmVpJPilv6dtn8opqIdhT48RP3
ynzuoA+R2yx/BD6mjyeYfGq6RbUI3ofITrAAtAhz1V1qPMfoXnFl8VZoVrq71Jg+xu94T+XuKW9u
5aGA7//tleJJCBBLQcknqPAzJKTE4GVNXZpctYLd0YMQP80FwAplQhhimPERJLbIC0yEEL+RBdi0
ouaJDPdYhK3QbhpNyB0kTAQufvVNDtpP9sDutRYIPSTVG2YOAzjzqpTnIKt9InMbXKJCfN3P8cau
sxyq3mkIOhNeWW3mP4WUsH29FfiXsh4GuLWmhP+UiM+L3JBfnJYcztzHOgfYJiCgQxKMSzfW6Zkx
zmd5Ri8ilVXJ5rxAmxSzT3vDMUzx3qPyU9m0fOAtyOJ5Phk7CV4lQXMwCh+uqy9DmQpHXwENr/7u
8CBzeWnV64Z/YwDBnx7i2Qn7aiFfYdlypp4s0Ziy7bQylvPQZXz190+gxQ38M2cC20N5f8s0aKDx
+C7AtuH9/1qe056x3XyLC+W8HnKGvEDpzz3vuInM87JmeAF7lG9V71bHHzYLR4b50tu5GfjiumXG
HeoWIoh1eVVLnErqAzJXf6E+MBJPHAO29GFlKU9/cpiUzTCLqSaxcPJQOnGfA1LRFlS4aYCy/nSL
q+8F5x0nOPPY8iDe1lSA3h6ZCisVUZSZNbjITIIQg7/QiomLH7bRV7gj34mZDiS2gx2/s2+qCqnX
SKEgi/Mr80Ac1Ho1B0DMIj5Hosiuhw2BOpa3PzG2xMNCR7IZl+NUimPxuCq2fbi3Zxfz5ermXGBg
9LVtmoQApjRdkHRpcbFWmfv+eTPPGNLjNFLvg5P0NUL5FRyer9zsKxGsZoCSRPe89Qun2BS+o30J
zHziX+4pjT5sXG4DEunXLcAORJMK4IcnHFz14tXOb42b3+8VXjwnjlqux69aGdwYmAbTrA1rPhRg
E1yAyEMgHUt+TALiisusuM1Fw/0ZsoboJzPh5wLHU8igL08YrdAh5fT6zGyfmvrUxvFlMQwCr5qA
wgHzTNU5AfT9MwmOpoYPvVNYuhe35wF0LgLcqwhIar7djaNqc7NmoUZbuhRry8M3jEphbHjgQL/V
JWj3243PxvR65pB4N53Ec+C4pcZhp+t3MUK4+ifIVLpX4O2OShWn4SGFjtbKFY+e5TYYDiM1mstL
uv2lJ2aEdo/EM+iKZmWxDbTytv6Uzc2Rc4HAyBwFHg+paAEvfHNMCb0K+lng561EpOhrVACy4FSU
CUtojIcfYg8MZz9xWK2iSrRIloTYPkSfNirClJyiDMZ0KlsmMh+ypclXNK+oVoSn1WbbQiqroS+8
C8p43vuTM08CKmB2s1vQjCPk2wenF8jx/zJKd0bd9+t38yz/GZI700f4DObHC/2TMH5J7wvfC8QO
aMd6zsMHWEhNPBy6stMuQPmDgEYwxVi+j8hFV4oGGLmo7BaupoSe2jOhHIxT41fGBoGJPDDg6xDj
YTEquCDougDGUg0FNLCCNnFNpH6ok0YZ2aTgx7qPHPbYsVRmLWVQzQ2IxKk7NMNbBPLP3CIXnTod
vcmkAVO4RIlx5bpT+7pxaGyM5uqNDjHQrs8xjgpaPiNrBSywbWemi9pH4ATlnHN18vKNSvUbWr3u
+eJbuSDW4gh8SZLw6UBQ+n+8y55gR32+MaMjI539nwV2QZkFJ+oPOEI4sjw41Vw8uPq+DXDqdLjW
by5EcXA5kolHpWHq4YoWmaOH6CPIanSw1nCaKb61X7WvlJoEqgB99hGVGZuX+VcNgJRPahRv+oPO
Q1WvDoPaljWY6PelzQnIt38cAhDTA85JsthnzcwcHxuN0kWB+u6lnkZqCz97f8m0ZeA4rwyARCBE
yokL/igm9TW4+O7PkGbet41fYojAiDLqJ5WdfiZjeJolAPVvuj2OqCMqr4O+uJehH9fqWNHRQeuB
EpgKvA+1pfs05HPeV0tUJ741KM+TL2wiQzSQfTSt5YKzwmW0eg3tiUvQQqYQ9ZtVOq65tbb/1zu9
kR13hKcF8NFe52ODMNhD5iMnuY2IVwVOIOgMP6Fy1SFC/s7CE8IHWrPCy35QbwXfhMj8Le2QfPtw
kUzWHkU8XySOPSWdcgMqDL35kxQdbuvAmO2JccQFw6R3YHoFgjq6u7+uQVdpEmfc3Rls/DtWEC6c
IAtbQg3zGKV2NRYWJZSbmo5uLZi2qtIOzly3e8geSot8ilv36HwPuGeqDSfWf8+rK+JAnn80Qc0y
OMrH4egxbL3An5P72HAWahO4A+NHYwNmkOAsy8sUHZe0+mdUWu4ZbkTnma4zTGLLG+rBCqYTpub2
M2TlMhKdlWqrQYYGsWk131x8lTV7+Q/d5NGqbgkMI0vkTVM5fLlEcNC8ylV+fe9wzFNju23e+byu
vluF2CpGO4N64ab4IcsRzWMU8o65I+DNsdKOrZigEOIemjK6tm6dqPaomvzDmlEflc5TmoSeKUno
PoMaKA23kvOZN+o6HL85Z6rF84DE/HlkM7o3M38O6lmxdyXixvFiKrTBe7brjWuagyKptLrDbbMB
dSu15BmwuEE7ev363Vi9DCzonaLdVveww/B30rMUhtkC84YZnADeExCQ9xe3d/Oe+E0pWpFkk3BT
wnJFbp1KzUnmIf3EJcmZIxB952epSuFTjsr8UWQVQY/gOj6CZhcZJbAwmSPhSxOxpf/v4m+IVjmS
KNZYPQdWGndfK3Ec2sfwwxY0y/eWv0V2IoGANEvpgb14eCCYbyX/gwstq618bSp2jRXeboDoYTjB
NyomwdouQKZLUGPedaUCoDyQR09cCkpGT0LcayzqWdxQ/IBy+Dnfc2kyOVraf3zXNi9bTLaNg2dk
JRuyQ5vwxgFrKZzQeDgrsdg7eDvtp1ocpb8sx+cn8JOM96Qgv1krlfdzmQHoAg2VxBi4udVfzJ+l
lIMF5RLVjcU/tSkTqd8gJu9y4SWDX2FWOYQyR+vjmJg2J9Zr7dYtu3Ci1nrmZ37zVDmuXQFNCrBg
ZbCpP2ocS6PCo8cJU37XuYKxEn7+1POqvjysU8asXG+wHYrjBnPLjEtw9K5sFpEoz9DlfDe2sQpb
c3zh8O761enPSbdJi9LrNrTti5qM8glSxUCdcmUwBDh/LLiTnm/mX6vo/nz2Cbe3V80saMrYOQMO
VG9VKnyGHMy6AOhRxY+mq7gKCtp+FMIxEQVtnjbeSxzbJNxgt/7slCiyARFlPBt7U/dJSTr1UIsq
1D6++BoOMmAXZxP5oq5PKTT9AUtooU+uvGFnCwbslcpsf/SyN7Hahsfga373c4uozvbmOUkTbAo+
fPM1bu9WlcoX81kRo8lQUnkwuDLup+eTgYmHa4d8BAYUjR2agG0dIfMfXtVmsTTzeHCg7RapXYoH
S61+mxGGfKiGHsGyHfr/BG/ahg4r5bQLXNVIJdVt3BiHnRWQlJMkKWTAGOBtQ96a/Oc7S+7htaAE
hzj61vDdXDTwj3IB9xjKTSuwZnReygYLbCloOwKDGCXaYuIedXLiqhuY4y98e5/IeVeq9k/RMmV0
z3NlOSBzltne2RHztUsmmucmSBteYSgwjdK8etmq+53Jv9K/Z51+iAXJjEMnxUtrvQlJDANCjZMg
IlFbPsZ4bVGQE+bXvLH94d8Crvd1JE1Vm1dhffb4j4FatU2F9zktGVrtU58H0xlOoT4nv4TFUdz+
JJ318dFsz0MiBNqIR/bJZTA94oSo6CYzCzBPHCQDKvA+nSesVJ5eZs6gMEHT+q7EVtH6NA9+kVAl
bMMgx5ksga5lTHLARHjXRXz+Fn4qdIMyJ6MpoJhVBwFKagRtduF1EkLc5yZle5WyrYSYZ3OP4h8j
zxlv1JNen7khADlkGJ9LbzOp0in30ExW9sj3Uk11C6xeomCk0S+L5zVcvFFhrpnAayl77HaJDcLU
SLH+9PF9mPHNOWL74VpCQ9t6m5y6R3lVUifo03zvBj5Gtj41erRv5AWe8/hehHNxbTTEOCPYLfOC
jh3iLdXOIwVbSbPsRZnFxt/fiKi7fbCYT46j2J+5RH6WJneosXhSMfppiMm1/XFz7RYDzroyPO1p
9ngV5ErM+nqQmacmnEGkwPQy7zj9qT/BM6uw38pkJ3YnNq8ayuafIhO7VZzfBAHeEITpRf+XZKgY
5b8IdIHGIBDVkNXs65wyZ0tmx6Dl0I5pv4zNj4cQhNs4yBNildl+OKEEat4bD3dAo+qASW6kvhwy
rO94cdeBdMeSbPGGy7lCaxx2yOZK1c+jvfr84qIDBXsjsybjCu/j7s5ZGBV1XJ9bpW0Sk+SStlew
2rb3WkB84mnNRDr/E4ePSVOo3Fy9AKb4A3AQ0loWK4KHl/tfhtNALyoalAAAhLgi1VhI6UKaVAjq
2HT6rSJEh5BxS73zMlUW/far+xVhRECknTyLWCRhn8v22RveV5OZ3hLdBjZRBIsx2lQGn7DmS/lv
CVgBAeNrat3q2lMvy6rrHnZahZERP/MtFZVT+1N1ThUtFdVVWSAAlC6EwSaqeSnrGKphz/NhwfCF
uQ/EGClM/t7M09AauhTyL8sjElCrL4w4zy0Us1guhIZWQTU++obdCBluCfkFM4yN1hACwiM7enRz
EzJmx7XM3B0s9MqI1v1PmMrGlY/ETy5BmMVDowYu/GCw4bg5yhVQozDG+pvTlY257RMlCRIx1Ofz
b+Apv2Y1hzt+xGQPK0GkM8xviI/WR545J8rBaEe+G2LsHuJ1U+yTjm/dS/if8qTc+z9HedSlSAa8
eoihKDbylXYOY02c/WTTk0rr8UCZ5RO3EKh31yjyigDxoJKVbM3YAjx+vv1a/xlo6XqA3jGKuFAS
uinsiq/zDPVLe8RciFgLi128yLlDTJIVa1wlSQMlUE6Ca/YWZDQg4bVGJJMFKcD3R0itsSeChzxE
1GpbfUXKwQdkXetT9P4axYggDf9KI509h3Qvs//34I3aMcUyO+UcAOmB8dBxd8jCsHLcAiWRBOZA
WHHyXgGL0oomyPssSmwmiGT8tZ5W2Em9KRiL3PJb8xk5XBTtVU8ic2etmScmKQFuwCElKqfSYY1L
Qy5wu+DWdC34KoQD4AATM2vGiCgzsTg+wZ71NxkZzGBWueadX8Xkbh4RXzAs1mAYUPdPCZOk7q8v
pG1gIOCXO/ZI9BcfPIUjNVDKHEfx2X80P7ruBx5OXThgl4Nn8U0fNotj7+9IsLYt9T7BUydhZc9t
ZRYy+QrYlulNazuUQvKx+lvvgcFSqROerhJXdetS8ZSJ04SZsyuR5LqNm7MLR6heoUR3dNWsloOG
A55FASi2HGhfQVWoLuVJ53Xf8122ex+qsDGWTvtgWmRDWPEeIZAb70wbekn51LGBpoAHPm70hVVl
tkbuzYQcPY+AL0KIcenddHyNpSwi6fGV9AjDmHaQv93NnT5T1IsLO0SBVKDyqtCI31Q3Z9x72a8g
vDV4aM9NFDPEvuy1ir6jzUdc0nGcGh9zVvfIbMupWL3mNVbHTbCbJUh1dubbjgtvlvIjM+bSBVrj
YAzAL0KMwWas28vcU+LqeIIN/Qce0M+T0L2A7bp240S/xiXbXI1681a0G1Muhc8xP++Y9ZQbEx7W
4HKEWg6Pyly366Au2rvwFWYyi8pzL7dxtv6VPKz+BBFsPy7kt/27NIvbkkDdZ94O0vUXAy/UJ3W5
dd8L8tOOAm9r6W2pHnbpZd9GIn1jOa5wY2ps4J5HC1TMr75btuVkEe/IeqY2Xlul/MWqLcnfqFcC
R+l8xsRy9VZKCWtKFqg09DPbfzYwI/zYodpaBVEBU2HTbVWPjmqHCtXxJ203mVeqWtHh5HNWfO9j
WR+DG4mFxnrh2ewFuzbtzkF4AKRToZatIr8Z7MT0jdf0SKO4vXAe+heuPPujJVJPTo9FfGw2gapp
we0MOnwkrWLKc2LROejnmsvwKXjGXO3gt9ywk65BI1KBwa1N6Hxs0TCNkHu8O0mQETi5c1KF1+x/
Cj1exmBSC1t9LI4+Y0bpHBEqzFpN+lo0t59imPOtvmxPsBGKKi5WFXClrZfqDXXHUd3cUuNS0eK3
UHEr5ZC29zTh/bJZKPi54nYK27fGs4lejcOw9sF+SDfjKO/IUCvi7F00rMkDeW8Qasgi5Vbr8RlX
zW8r/GLNoD413VCtZiGgPovYpEMEhrBcbt2fPasoLPgV81Y3OamR84Hm6GYU6uht3zY6LBvfhK2U
LFesB5GIeD7Q894+POBqXKGnsfgU/C6d8277N7XkxSF/tIeb0AfBk8Q00RAUPbiX+tYYpzxWchbE
tKcswX12VmsGU1IekLk+ydfb7+FD8mSif0KdeTRZTpFpqu91K2tkz+0r6qhU3BmS1jzd8U5BSP/t
T7xUe2xFD8S2V17EAb4o6MCDA4cxugkIaexlZpqvyNiV+3paaTfClVjbiAvo3MLp6qA5kITP8u/j
Oh9vkUykgbrQd8DxqReKJ7l6eRpA8LMTh4APM3VP3hzlK1ddm7JB0mmIaQodLwGD1w6SGzc9/Jsy
H1+LypTgKu4D1PS6zfymmnMkJbP44a1ALMxFtt/z0mlUDR5efTKK9XMEGLdfK7ph8KrZ1m3V8+F5
Q8V5JAotNqBZZvHzzHWJ8wUS5SdLIftwqFA8Be+Olbp7SPa590fRmQSnvF8SQRb/iuUdHgPzOuzc
pQPElzb5a29WI5Sz56EsfdH+LkNXC1zcSlsE99rPM6Nsvg28bG+M39Lgw1IEhEVXbTifXZBozF4w
cHYpm6d/rryOtDodDYoofpS4MavachSdj52K8yIOvdO6Ma3tdeuxD3rmZEmXRWfMQcvVBAoZudg2
i/qB7pUE7+PQ5da/qUHzlGERGu3PPb7GE31rayJ5IfJz51Vx+z8lLRVQnZVI8kYsFmX70UEyWPf2
nuTG0xFPbLKs4L7THoAzPKuCJxM0fhyohM0uVkY0nCr4rv06ZPMQhPpQ7pzYFepI9O/5e23ezi/Z
vBI0hCpC7HcSQwJcmkHnu9kH9PtyHSNU6nsL/8oMZWYRjyixKVeYYB1wIMCVdjSPIoWd2LsyiH6X
/++nUqvyyGspjGm0Ngtgnrvpbzs+6pZIDdEY0bB2Pu7/a9BhsCjy7bpHRmHnqR1BKzNP5YCxjwmL
JgidZ7bv6nEKd7AO3+zOuIKP0n/QyrfG7SJmNbbCUmyH96V0OimZSJLpElfhGIC5NiDTfnJyL7Sm
pJBaI3GZRZYfpTn9hkwVhl8KtnC+MCfTng61uUy2hMhSYeZKCsH/doS/dIM3S98kdKOEaAqy/XEm
+vhFcOp9OFQkhC/GhgM/mEa4yZbQzjX49F1jo1YHh6ScMDuzw26abDd6oac/L/zEkKoXF39V8EwS
1yaahDCkMbaHSnWcatfBkGjRr42U6ciJP/dIFEf3cMLMBpmzD3mnxVswy7OhTuEv8P60HaxdqXGr
XRSVQrzNZLUQ8EJxzqHGIWhtvtkNI0SAQhMNtN2NMkWIytTJjWiCAAyVz27xBpcmF9A1p+XeDl9E
5Wg1Ol+XUZcAR0dUq9Je3ylXOmq1Vl9jA8oK+Wr1/Pd4tlHNPF0l/zfQLgGflWRd/4ZBaKA5Bbrb
QZEIcwW8p7fHDJ74aR+G6JF0UT91JkdFyaqoU1wr6e52QinxiQYH0xJZlybKjb/XbazejdNjNc5e
dqlkdaKU+P++PONoyk0plyftfd2KTioQF1k2pIhw6mZ0/oBUzLP31F8yifm5Pq8DBNzJulOJDCQQ
vC2PadqQt1tbSIXUAO4h8qKKt+67ghOf1idfF5Z2BFdLOe1evLblOlgonzZ1HSlbZL75KTcMAwr3
iV0OQwmWcBlG3NVsJomBG7VKJmlmkfJ9wHIPSALDhcP1FXKSdHq3eEZE4pl+EX4amVmQtPbYei5q
Tll1bC4Abcvx8nUki40cnBeNF1PavydKsjfAdhBPS3vGuYw1729ujCP8ZR+GAAArwiHyx+k42Dwi
63zuAYPiNzdCSyNfABO5pn7kI1aqW271PQqn2wjwOioJSzM+GJOBe78m2oVRLtJuH+/iCM3r4UtL
yIcnFbPtxO9lj8siuxBqW/cg8D00FibDFmQmZTyEdJ0hGP2zrY/oTu9XX3JbDEwG1CTKTuxvM59V
efOgNfH/nCdwkVUWDUc/7ILIYE0JP1wLvfD+ylq6XKuhLsvag99JEsNwb7ufL0SwlK7S1KgrTQlm
tlvaV/953uf90m8ihXMxk1Xv3+/xU3RfnmVorig3TurhL4RdWVqy2YPLEeeyWtFBbFOR8jeuUcnE
ntfFDpaoaBkWIv141jGZbwq8uqiS7ZazZHaC+pfX7GYNDmMRkIwkr+wribBZZABwt+j/OcEacl8+
MI6fOqq9jPKedlJ/7g9ohCmyBQyuW4gQNrnMdFdq9Tu392J0WIiK/NRdpgUk1NPqFRBQKgFBrx2Q
x4XzH9jzOY2gWGlT4zZHykwB4grpX/BOI+gNu3KgNTHYEKo1fXMqy6tfy7ZIIclJd/FNZJZEZfDF
rvJ/Lv9JHUAsT6aawXIZYSknguPyqXdIvu+rh2+3jZ9U4/WHoMx91SZhEzxLhElxSVfqIQjG4BWD
q8FbXanHVVZ0FsuEl2XmUGPcd7ajdQ+OaWjmBbDJkC09H0CBN463hxluN68ZOcUkl6z10lK80sfS
ytuZsnOi00XKARWcMgq5loLxVFdpFfdJhhz+7exmCxlze0iiLqTifN5ANz9p7YOOr4TEcjwaTR0N
miaAIG+eJmeCd5sts+JzPozf0AECduZ09jgZHACRXExbJ6HVmaiWgrzK85yd4Sb9VWnKN8d1if7M
p1tGBPGy5rdCzMtcdhgvz6RsAsuIc3GKWF92LoeUvRN+eO2nKJFk723VTZ/vJca9/j8RBH9k5tNO
dQFM+vBOsRtXA2lVsG5feM/AuLINZcaz6fxobXU4QM8QEGQZQYba6E+jL7dZMF/7BTjDhA5IQOh5
iCk6SXy+JUa4P/IBDsnE9Aw7neaNG6O7c/lPo7Dr+4LSHQxbKr7zcf1M6MDQFEk4S3rtgCcY38Lb
ieOoiIIvt6Wgkb5c2s5PwWyuTJujEzqvQ/yA7Foiwbz4Lvh7lxYaY4Pfx7GSFGYyL41K89Q8npkQ
WfZTepfrySVcQQ8w8i+1+d9lq4Q55GRSjkJgPV8V0jujYr7Re3D3Lc6WrI+UU3CJKjnbgZHYzGaP
yEEEcy4o+1fScw5prrl0SwtU1dOwq+q1QHF9deK2mRliFP2oM+qbRk1FLe0PTn9Qz2vAqvYeQprx
XS6BqRmtgYYN1AS1S6xmNbomAFe+BJRBO6blZ7ZWjD6thkSWroSgTnaNwHmIp99asKh1m61bSa2S
8HA2xOofoWvImjtqq0ZtpZlnA7mRDVlhgQsr9NDk2PThb3RLujn3v+U7Kq7FvJPMi80nrJwng2K5
ZoYhXAcoeV4UmoZKQwDwOsfpVJgRvWhC6deIgJhsI8n6+oHWHZfz9jD7k2UymgPxoY8tPng3f7hu
dzJId2aUW6fVhRfBtfmUTD3ycC4Tmls4WxsbZUKizEIifoiakj1uZ3e34IuK2cvFfsRLGpcW8ZDz
KrlFW0xHvIJZLguSe4HwDEMoN28uF890BzwnGDDNCfhOC2C5oKwnoc2ArucqT3SGgJqgIThUc2nN
4PBSZa1PbFgvI4Ioyw2WCbr/61mCNfEarFMqZ4FPVE4lRQM321tqxEhOeFlEIyxR9YYwUq9bljbH
11os7l6Q42WD3ZazAjLTsigaoyg4W+2rATWay6+JBJKicQ0lRTTjo/CmrEkZObOldne7A1ImqZXp
hmDVXPQJCocJDvkwHrAtIAdJaZtwQ8YYSouz9SYFuBMOIkVRyY/KbQEUKzsNOa7joyh2ecGY6A5G
PrUHrXZ699qlQyysuLpdu8UJcxgW/TzPgxEWrbLq4kxn0zQEJ6lLId/B61vZGuf2As4H0xXkpFn4
N4KVkofpAAyaaNSAXPUOvSt1btPuJOOntYjKYJ5iIHdNjirbqce81dHJn+UpncWDq+GzOpDDY4Rd
2WcSEeZ/A3469be7spYDUSUQmtaV3aC1Lv8zsgDhhdAtu/IeDOK7WPCej8iSH0vOIyVqEapkoNF3
pGbdrP65vi5KWvyxqwFald7Pg4gmCGdKoqCIuYYkdclJsVCFqcsF1fNH8EWCWw7UUaNCw+YKKAkf
6am8HuY91sNsT2ztSdvROq7fXtwjnxK2eGKkq+rc9Qqq5b2RLhxdv+WfnWNf/jnmHMV7DHes/GAR
LfrjoH7S5c3LHYuhnnlQITYUPVPWtCEYHKiV47JFGc8uW515i+fpXGwN6E46Sen7Top3gpa7pD7/
MdCOjQrbd/yOrITMFpmrvrgPkMZHy3FYQ8LHDyI78tj2NVxNjl+jduFWS9B7xbbXtOn6JEeQpHli
FHOVs7CVK32y2MHw7v7I2HpPYoUlcB1NRsKP0AF5Z4zWh1Q6t1KjhJIOZaz9gmcokD1jpjz1aHvA
kR84SvlP5hDxEsR5BxcPurexILMTWDUdohFXDHV65l/idiUgkDV+IHeOPEACFSr4d1Bleqp31duh
Dib/kEN8hWx+mKNy7rWkyU+6oREaKirG2SK2dSH5/Kg2ogjRlomuRKZasfxaCUgsTG/iSwPWpnch
SXuTgp3eiVSqyOfVr8fQs86j68o4LPcOgYYeAO30RRi0sLImOsJe5gu784egkNKHS4cp6+QqFH/l
tACQDJZMsXPh+Z6I50E3RZB+jqwKAcAoQIJ9Ns4wnBUmUrK+DUK2+lawWzTXt3QD2zWePsb1mk7o
5J/rmZbjSn3OCj69bjPLfHnWYCmNKhBkXVTqp7hBWmUcXpO0ZDeU/u78EIay/IvDywctEs41hzD8
aWeBx/o5r/Xa3tRVAfrcXpoPxm5dRwr8GvCXNwZmFq1ZEhCVciytnKKXDmD+S26uortq8m4qcAQq
ET0TMTqRqEOu+NIW2hUEiiuZfoiFAePFBemYRs06n+l36o7xxS/pW6i+AT615jcfVjSs4uRuntIv
9rvytbK1sNjLGjSzTi0IxCMdPK33mSUsGSlKx1CEpUtSVmpdFcjc06SuCviK7aaTVJ+rZNBnsSvF
sTR4Caigk5bMie0zPc4xzKe1x7kpjuEMQZo0NWAwvvcfMlc8tpzTd1h2+qd40sJvMAIU4ZOPjKie
yJxgbW+hjYtfiwsV7hAXWATAZfK66cIPsYkpqgOcIKEudBEyPLUWKHaFt+XOX5Lp+6lD+89EYEoS
igG21m8qK3jAMnYe2d7+50OI1x0afoONfbK1AD22FvR4+G/7gTqUp4z+hkhD9Sy0654Mt0rRwjcu
JAASutsQR+Ed6GTDmygv1YEqeHNpZpYn/Tj+jK8iHXuqtQLW/yQIKB3OhvojiHv1HjYjA/ieQxrr
uSOUe2agzW1w3R9pdbJ3OdQ8LmJ+6M2Gw81xa9veAf+ATAZNnzWZw49NyrVLBMq7M8fq/0rvGpPE
2RGvc9NJGWoyj/6ETSwlcQopfETr6keefAhEc64+UvsJv+vZgQtpqrbCXL0OPK+biBbdFFqr4S19
tu6s7c9kk126vt23Y0KccxJx+yNOmnRaop7vWDcKsnFQxYXwUd44HLIMATOj64iMi6bPj7n7Igbp
ORq8Tt5W00JgWOfxoBamY1RdDrFPUY8AAvASXZmQu0nMGksMNpfNsZdLcIjeUcIcQnnMB5omNDNF
a6l8/xSeOV4g2P+IM4uk8QWCK2XX8DqzQdyyNCKM1ULR3QGQ6keR4uo+hZ6fjhzFmlZWirSqJJed
wCqrzMSvxsnlpqOFxI9FgTInWfQRX1u/4TX58RFC+E6FLkgnQLb+QRiQFEurQ0v6pSEL3KJJbuB5
/OiD8SC6xyubzP2U4yAGKqpjxnIha3Z9wnlppWryBA+Mky2NEquBCeSxPSBFotJv8etN7Qv7VGSQ
v339+cgeNFfx1EL7MKmk6eRaDnF8UC6cepeyPAPZdjEcpYGk4Jl+LIGaoSJPDCBkdZuHW8uplsO+
bDpzTmG+cy2n6SzVEK/VPpEK5HSCEzq3Qt2I6OxHG8KbS4WeHLeoDzNn4K1Ta8M6JTA8RssvSUEG
n7utdAGgrXkivbNwHE/Bp5VFDZ1gXouAcsgr5sV2iGffnZKHKQOA9ZVzeF7vBIUhmFzRijH7zTZ4
cFNaMusxhuZxibt1uAapnQC4vEJQle6BwecKoODkUYN3Byj0ia7G2Jh52zP+zFLWkAx8nQQPA2D9
Ch/tehSj2DZRPBSYb1Kj7P3NRgTHB9WntDwjrEZ6YIGOUTFzyrB0KpYu+R4LuHEiZTk2X9QWL+ms
JM/obPzDEdJnQt7CAt+9mHGalGZ0aaFvK+0wciEJ5JOcVnshvy73qKhr810hNHHVEWVDp57XLgXv
NTp7An+vqAstzZ5+5uvmY+VI59GspfFv9X+tho5e9dF3/juFM2VEDQ+tefHRj3AxAIaKb4akzKO3
9L2bfaDpS8ce+LekengO4VXpEuJsu5SjfaR3EB2F2IVxxYHGCJsObHQjSR4Ppgh81UplVUC92iHB
b6AZAV2xSgPyvDwXoWl4h4NelWA2KjaZmADKeYH/DaLMFaEaDIW7P1pyuMG5ddNs9EhxbPcwMQVF
r73kRG4seTd8UAynKM/Jfs1nvSN65joBmL6ff8tOj91Eytu/1zxcUwl6Gn3i6zw8I09FMgnOLzeP
qwAh0VBHddFItuH1njHdTKk89IEG88S1d68JKRkQbBD8WQVdTvLom6eU6ZBBATJPOLwzfsRZ9YGR
cYVwFfHQpFl2qpIexZOW0FPYVVwWO+brH4hXVRbkQYq/nn1HFFSEtqDMA/qooyaoEh34PU/0ISQE
Xj1FSdSU26Vhgnj4PKwqUWQNYzI1EkedzsFL9cGz+TZ2ZzMiSv/f/r2sYTerDNk3OFsjrF2lTYU7
ST3k0FUpbVkP7pCVTUm1ohWi+ZLhw3PLqPVLaK3HmyJhYSx0OjUhuDLL0+xFIzQNF6c3CeRs95Zi
tWP1PDLWkwgMAYSWqoQpao+YTxopf/4NQSrD24N1arRONIiZNxaEEoJQV6ti/0poEguPCU+RhZtt
l2qFQtFmhLvtKn1Z9/6zsx09iTDvmPV92xF6KUmWjxWy8TyR50NmwAs8V5eyMxLpGGY2edoS/nAs
BAgH7hDg1tXPRMxMm5m5NiuGFnNIWZpUUC35CGAsw6s8ukddPqKS5YSW3WgmGiVS7sifXqIMmSRf
9lkQYngiz+ZRqYIRhdnmJo2OUSjX2bwJOfatSlWepzrn+vPBCDBMYhik7G3DqKfjW8YC6zkHPaLd
XOt+fzd2OionjKn8gflJbArjXcXRe1rXiPmUWBHZm//p24Z30ZTba4LCGwW/az3kk+TMoeW5y5SB
UFThoR6+2fQWgXEBBO7xvxk7yiwX6fAzvWB+3eSsmnF3hFJ7h3InqmKbvYHzb8LY+RZbN2vM/aCA
/nBKcfHzij50L9/nsUcLAmylbIabAGa2Ibuzwh99GZpGze+perSGQlNxEwnzIUcyc59Tk21Lheqi
pcG8ggQT5h69gkCrA2z/EVaOlFxrVQ4uAGZxjlXN7nIsUONZ+lWOVtqKArCP//W7OORhbAbRY0X8
F8TVVqQ0DNcnwsA89Nx/m5uMYVNU5MHtL88ipYkRF3SPWgVz7QyiLQAy7lGq/sk3AP8cVlxUU9in
b8P4WzQQ3oYtR7+MkCi5viAso61dxslGLknkqPSmZkoqJSp16IosgKBo1jsham+WZIYqnd+Z2Rc1
JxcEwf6egooNRn2alm+dF4zYhdSMHKVTaHoR5lthH/zfh7Nu5v/7e8HXSggcUpDI5Vax4vGdG3Ed
WIsMnj2sweoig63AWcbktOZDOD5/9361H9w2VN6ZHZItvdgLXZGYYuvHcVy4KAO2yz8A/Hhkz955
Y7yzWEZn0KCW/ld602brBWyejFpQh/J+XXTRKwElrBIS7kM74kWVTJoI0geKvjAXnrHhU3goaqYc
FgCGTYXe9FEdgLEKB9cLUX9JEK3RbGXhuQL5nZfOP+JLHVWq7bvhWbfab8aGb0O5c4jWL7PiPcyW
X7oO9RRMgsFBUPnTjswIqPQ/i0nXvoc3uJ8w6RMYNlU/GWM/0HghRZLUrx5v0bP6Oem+fjuj8yIt
KyVjHg7QVhnc7+UVrfhErDntJ1JMJiUNn01rZOS6EQj+PZE8b43s9vyoRXlIIxuT7x2533ookiHw
g3Gqrttm9TGUZNL2iJzkAVLVSW5xfG37+GiXpU2p47oT7lHeF7ETpYISHJuIZWGHyonwGHHTssVg
jaa55zLRi89PYZsE77DE5Rlj7KIOjRh9RxI4NC/CjNdUPGFB+r0OjJ6EWl6D7WlK5uM0tnSHT3K+
Ro96r7BkJV8dZiPGUW5Hm4MV2MBCet+h+EibX/BldR+SLSzj5pUlqtPIVc+049mfFQRuSbDrWlDe
brCHI129wkHHxZzlF0UITRvqJq0YSnV+QHl5QJ8HJN38nEuFuOq0JQekW2CEkq9ZxV0iiK5GqiPc
Jffl1qbPR43KjD3Z5/oDuos2Z0j3A+RpaFe2x/VUaHete+ip2GK4tuaArLj75uBaefxQO5/5UQPD
AkqrIsWmV/q7Jrpi7hMH6aUheBSigI6AGyOwcejU6eON1RfaCYxLh6gFhAhmiqfgepYgW8fWcexY
NwzR6pCh4vC2i3QUe5HW/em2PnKsiuDxJVTF7rC5DJ9mmPMy1YexPUoPUzFxq+fJcvLbN2yaVqJv
tvsMIpvEAogSDPbgzcYISINoobJM305EUPJlPn1NrFVQzEjyCWWPnzx0XIQtixpDMBTzB3ACeWGo
XqT87BwSthlygKMFprrWNri+2cBlfHul2q/DxabxaMEz8LB1b72ZSoHAnPZdZD59KdL9kppEl3sV
2OExiX2fruexbgLtf85Xqtr0jkWcPfWO5nUXN+X/U5Ic5V5qQgGNfGQEF4YmJ8Ly/yHzNTE8JKek
HUzXg92G9J45qODv9FYohLdWTKLRLFdlc3Hh9F2N+byVuJhGrzp5XzNwCzxtednLdbzGCEFHS0mG
JFc3RQdmhSAlEWqSZ+83edwzkNQs95cO7Kjya9Om6cTnpSu7St4d/2MG7KglAuJnxkWF4TgaQ4L4
j9JU2G6rW90DfS/uaxPh9FFdmNDzh+8TXGtLJNsuYwFWC7mfy1s/5yUqO/AF0hdiudq4LD++wtM1
21YZekKwwnYiooJrqbgrh8tWq1RzsGZR/LaKeXWVt/m9yLg3VBna3e2DisAoiNgQPXmuJBwDpZD8
6PQfnvLUzfe/o5EB1SkcyHAjhB+wAcMSIdYd58Il/jPn0KcF2vz6PV/FZFe9vbmZF/27cRVSi3+J
Ita3JJJEWwpsJGm1hWljIe9u2CTtMXKhEAilAvBk7ZIvf4ujMoxiRBHb3eCq2vye2Woxy2T0z+0l
2R+IeqGk+xgOkh7UZap/GNL7CXL0YW0qhyc8t2O6LjHwQwpqbBjcBfpDHMDmlx7gGm0qDkQ/WQ73
VN1h5M2zh/haFT7+cNW/Hihn5wuSktAzH3P9WRA/eJZR/LakoUPCb6wfxpBiIBbYNVkWrvUspT8p
jYYYoWP8/yZ13zrTf2zHBr3ZgnY8yPsYoMajQc4GqUC4NmNs7/0A0vnpvOVcRPx/xVxvrFn0aF+I
MGQn5uEGBvwRi/xhrsiX6c68/95cdPC/CJLQ+lS0HvcjGCcZbgKFwSnGGt1M/sxMsDiFo+zVQI6d
DW4BTdqbWrePp3sOZhByRmyiQ/RJNF9OWX0ymwW9vZx4R4al7ahzU8TQfCbY34Yv8fYqhmnV+1u8
2wdiSmLLlKMbgy1+YKmE+rh0MBuiw84jUbdFsggFSwg5HZf5OX4ISdPULAAs05F6ASKjNWxJnB0J
V3Qn9QljRlnbviR6Fj0ak2TOyOS1LLZxWF7Pzy8fcKleIYXKrimgoMUwNqH+AdJStqjRFYLVoxPt
CV+/yscXUaNamUDs6vjzHUEWjZqjeYRauWKd0u1mI58/Gs7cHV3YfjZjRDhY0Kuo+0PtIY98m97K
CL/NZWax7XRFGRnBQYWt/BK/P1cvaH6UujfnEEe9amMHcOX6Gcpbh2oHLzBECr9lywxb2XLb2I8p
xCnUIo+g6mX1T6Rab6cS2qxzJ63y7U+CKVoz7I+9rRTdHwDo9fr6eMi/aKRTsRWjDsOAQs+vjrVB
HrQKIkvDdAFkKphR2qSyTykrmokuB6lW31j9PhMkwU5i8R+oiAkvKDKUK+aDERQf+Lh6ma50qsCz
ieLes8Ac3p+Jh9j8i9kwCbPHPvQok099erKXxlcs0ouOuyYqRSHGS2HHC4m7bDq8eEEd6/2pGUVk
ISqeBdbf8MseLSTxi8i6PaXDJVH05T15CliF6Pkr+avOHD1EdVzpPYmvHH0vQpZyz4GBUiGS+Ux8
h88UBWMuSYlHkcMV0/V75gdgB6EP+d8zAerBNmx0YRgo7DjOIX+6oRiJ6EUXI4cU/jMeBxty6we9
k1X0iCj4JMGp0YuLlE7el88ISLsXz3Rd0Ykh3o1qrnjSi/efp9UTt3a2pWhLPX0BkoIxWYlqfngj
uSncxvf3J/ehMzErWFnoIu8Z16fZi6AWhIw/A6FhN3qeShjokQCGzEGJ5kFR3f/9JgaUwZ8X+QKm
fzZRlaNcM2vH20KDGybojKguXsn07o4B/UUA50aQB8VJqRMO/TgnghiwbRVgZWwAdoJXCg/NkI+y
2OnOcvSVcUCwFa/aaYzT+hk6O661EkNiIHWI1j+c+zwgQ1d0Ln5g4fyw004pjeENN4T4H+DaofPZ
Wchw24jDiKgu8/blJjgR2DP3I9AHOo0av1CJRwCoGdwrhX33s+EwnadAkzSYbkKrg9owevIPQdbt
G4v7MxyfwKlt+LcLJrWZVWOIdIdLWGhjcRFnLUVkj4iW7Q8JDsbR4UxM7eZ1nQnloaGgQNQa9RTY
Oqj1Vch7R4xuVq8rre3Bt+L0XXQpe342UdiLZq9esZIc6N2DZFnN1Zg90DFwp3j/rh47Pj+NzSpq
hZWoQZINf6Jr/VFWoA0pNtD12vTsoOi/wlHUNCmgshvyiis8e2nzVPKeQjc1+BEoHQzDJMsnAFu8
FXHqeLAhbzzMUkA+rxRu+4H/66ubgoPPICml5vLoM7Vm6xqpFXPZCrY9CupJN8okUaLKS7t+NAiN
7yVKlloZvQK0ASsVi3Q0i1vNOKiXmsR9EXheU2Dm7nXVxVp2D/uwbdi3u0NicVvXzxEhC5GOIb1d
8nEr2R24UG58Z+k/QAWnaVO085ep7SkJMrsXe4Bz30cItW8CVAodZ15imp4tl/DKnE+YSsv8orpt
mmfezkiKr4f6P4qx7MCcjuDsC9nl/4IUVDsfSNIJTv99LTyljV3MiCG7yPNBJBSLrpyycCbQpSjt
nfKZdr8UZ2iBDvRV/s1Ld/2Wjc6IlhtLCyJT31SSevJsHaSkINNqMBUGXqWmnkU+1FkbRqjJwhsw
22WaQqWtHWcUOKssfa52rHfsJ1mqv/3AcqCODaJuCdpLB0ugDnRZmA2gVYYT6VBpHn1aTIAdt4gg
UzgPAdm4/EH2HqwNRkUI5gztVhGb2auVvKccjHQYSamvcDEbI23i6jjRnMrke6cG31XEd7PEG7RY
ve/C5taY/tNkw3d6slP5gMwq6f20ZyP2KMHRV+NaPC+y+CS8ucgTseyxUhU3Dm+e0IvcT1TTZq7f
QmWWGq9WMNw4lnjslqb7gpo1qA4DPZ30tVW1ensgmYOGJCOs6DgRS8C3bLc73IdxxFa8Vz2Z13jD
+v7+H+CM89Ru8LzzzpsHQkab9Fk41UtK/QJZNbdvOWV9xe2wyV+1lqKVuAKsQ1CyllLw5WCkwArr
RVS5negSBYW2BVe7nS/BLuXEttvayBahvURlo0cH5y0WEkxB4d3Zl2fXUnawbT/Hw/LPYINjtzSl
wFMYwBj3YaQ64V2d/6KHrrGt11vWrtXscxFXnUoi3YaKLF6Tm9KyVPUQcFtHiTI+iW7Yrcv7+Qg4
nsfDBA+drV+0GjokD8Db0uLTry/6MWakG+4bSU2/q0uQig+aFFK/trj1SAmckU3okNKO1PAjlUpY
M9VaOR++U+RrutDGTSVwys2lpsSZo6DoaiI9dGfPrWzaU2rSqYCr+5XdO6fmGKyn9LN+0PC4scG2
JYwGABBIx2+Km1WlHbmczHguNfW8k2raWEz9DrYQdDJflv0GuY7WbPzAKU6rlnhqI6evQGNirgwK
NbbntQApYtVJ7JVeTT5IdABwCiZSwxt/nr8ThmqPnTtxvyGKaQu0LicSb0VHwyYviNqrVQjUl9Ye
XxGNWYkUmr4eLdwk7++7An0lWV/KbXKSMAw+ypNSERdXksBZQLSByA7a6+1dU5iO5MgUBiL9bo3W
5vRwPa3Pi1tiW9snNAijhegf7ME1t+G3h6yLnvfYj6Vu8pLU6lvEtI4n3xFrJUTG7fSR8W/zJ8EY
FYf5QPpq1fZhJQkSrqyqgIj0RXgByviolKToTsbBR8RTMdD+5J7ik9/YkcjqyAcYJ3NtOwVp5vgY
QCqPMcGRMw2Jpz2KRFD7p+vb1oJoIcpcwcI9CGB7Uq4bNUWK5vkVwt5McKvEx3XLyflvEjVXXEQL
E3mESP7D/XyJ65ybxTp9REhbBy+Aao5bP5vAX6zesiNSHM+jrLZMAHZZGxdXoU4S4IHmppQT4d9J
B/kn7sq5ZVyggzE0qX+uLASFdGouJ7oY9TKraYYOlYRhvwcSdWiogxk8Y3PJ+xSqpTyOQtY+D+QF
ObLh/PL2EOhaF7sp95Y+WshuUeEk1XlZmygyLSxH/4I00WUNZZEAkDFlA3GEc/2YdL+uhfu4p49S
rirqhE8I/Oa1OTWYHiUcBfPKHR0pKRiunJwPxrFm1qhFk9OaICUXHU2oArxfkwzm/hcX15FhNjDU
l11r0bzqwYYW+sVhLgbZ04LSKpPLJp2+G3MJYvkYIqT+B+Ad5SiKOwIs6yGo4KZ1E6+QKuqIc7RN
2qaSqJHyBXuwGPqQDn1MTreRwn0mI6NtcsPQoKAV9GyqOKxDUgIaACKASGkJ1ozUL6iEY1bsU6sB
0b+dzQBsKHeQ7WYC20iRhjxfPo4z1lCpeIxL5m7gBLcrUluN1ghCuAIBqVclxOoZ9viZegVCn3/L
+ij+2ApyK5sd/VNMlhYC3KtmGMEyoJ7qTYTErxhmUdUiFDQ7iLGpZb/cemiFOGu8QcWcPUJTyxiv
L20h6omtx5cPx9etMEhmJni0Ukt9F5r7bkgB8ZqIj8lvH7DwNGI3wP0T5mYc+8im6a0i0reOwYFO
6kPvObI7DJXVe4huPxXJdJVceVPWIL8Z9lGt2SZuXmxqvi668siOXsQ/2IB+MIwMR1ih9aaNVFoK
q7dIRrS8NxGKLqZM7iZhaCm3nfdeUccS6LMXE3a9qyejVDJXvigveyN7uOdKJkUYOlLWb8f8zAJC
JwDBV0ZDeLrCZl7MSp/DpEnKp9Wzwo8APql69UYiktYidcqvCpdltXiY5BJuevcsl12l40vuDn1+
J0O2lm7RFthOGFk5fY7/6hKR434fh6hE4kI62YBG85D2+PDNJ2y3yMwTyLN6ibk5HCK4n8ZpRGUF
lyldJyVV50nnnzyFVzHVZHlv7d3XLOTZnstN7BOdzefALikf7MK0H2DNX8JRgXRVX3l9O/gE1S2C
JpKziVLDCU0foS9z/fZoyEbapeQY3OTs8Ff6olbdyponlmuL0pCReNGQaW6iIu7oM3ovakVsWT1J
KTlcLx1cD3cqps7jR2LmWyPTujbtlkK8AGnTxl9Y7WmEHDXx0YaPK+C0koGGsSZJk6tZ9wl1KVsc
sxnD9ajsML9so+oHvu0L4myqaTowDK1DYtuKXOmq3ODs43XKZDdVxtireORwYje4hh8/Dg5iSbFl
vxv/C5vaw2GONU89ClGedPiRoq8amBazcXjKGl0uMqDkatBGm1mVux6JZo+jlSXDXFcAxLqJRLpu
6yDuewFNn/goXhF1LrQ9WemBz0bUWaZm6bKPuDzQTWeqV1YSloH3nfGi6xi1bUg0MvJ4F5OQ4qhK
N4tW4gEP10Z1MgezXPWDzi+ezUph6mvXJagFlJNzQP8zh6nNZTmI7Q33H1O8lk4irQ8/Mew4Mgyz
XwSTSSYcG/5AIwKm1t2gXavFvBrpBncdl9qXbz0EBKR78DlxwlOz9iSagpVuJugopVp/1+scJVyu
GAA0BQRPqNCP33HnhJkTAlxzQOMpE+poGxUUT2ByEX4TN0CZjGS61FviEm4N3EyEg3VEMi+K6G2r
uWIkNZsrrf46vg/CbFtWrLQAh6szKBaJwPYEeRQ82nNYxS904y6xTGTpVamEQbdlzfq/R4M6Fm0l
+Sz5quCBXpOciVuaNgWxA+XCk4DROp0zz7d8L1nf11NE9Wge/lMSJDW5L0T1FDk4BnfzykPOmXKx
z5J+mT/wGNKlJsh3ogoU3IAtLvx1w5eKHmu7HO4fUfqh10IrPmeRaQCuQGDadVV2t2VkVdt6cQ/I
zfqMrB5337km8eeKysxCGte97YgQasnV8U2jC6qu1rj7igkptE4Jq7viT+9jgrLCuzoKq+tRn8QT
NSihNJiFdCvqktAARFgHmyBM7GBy4s7/Jq/T3um72fTE4UwiLC6SjGR+MCpMjPge4riIUoBY5gTj
lrTI06kLZ+z+AHf5vV06Rre5X/jtR7KLDkDo0meFPMMAO2sWrAGXoOPKg7qZ1ndFpn8A0B51ye4t
EObx9OJ4jsWEJVl+fmJsgMs4DcDBmS1FVmvcIA4lVJIeYfAQqwdyicoySyxXHK3LvtweLtd8Ey3u
YUg+wdJTmPH2CJPvCezMti4dPo3aaey/cAl6RdiDs/yE5TOp0TESqPSF0CDFwDGB8t+bqmVfUloj
L/eDxFA+qNMAOkIg6mCVm0qTi+ZXTvwH03SSSUXBP9V8XcV6RyDprHdAoxrl/nGnI1fIEkgESn4i
V5UYRVsIF+NkJ2YMJWFehDWXYb3etEaBvRFBuRXETHL1CLF2upKGH2kCF4YahYxBjFlVdui3/LkV
zRWshA23uglhxel7mOTBOlR9gZnBxBph4Fp928Bo6/zp/cJvm3vAjhAZGbhiBk5jB6W6SSRetWaK
ckJMXj0WTEfDVbX6zzWiS7SG9fbjQ9oF3h/QnSdVQe4Z4AP0Ba9DQLaz8pQ2GYxiZFJmYGbh97IQ
Uq/LIn87GWt1s1uzgNrZ+D/Ep7SYr7t5v7Rvl5BL+VGeFNG7lFH7rZRH7V0r+cn+ROotWT7jketJ
ysNpLdjGy9IznB1oqs2HlImcBXXAf0CxKQlQl0bnKo6Ml6U0EcE+QxXBKOvjR4PJSHvBFx3IV9d/
AxtGALAI0jIgAR0ok7qlKoc2aFWgorvZscYqrh0869rQk2IGvbqNpXYa1N5F1Gq/pjdzJLqN9Z1v
7SdbRAu8BRFUyawjtLoaCLgc6qObP/lLHNUXuEThHyB7mbHWX/fhkG0yIRJtFjMH8+bGZfGs7tng
PrujIXo2+lDwpvbmNoNT+K9G4lzIs8USzZOmRYHlPYw997o7kd1vfMDTp65hIs3e6bzPGLFxkr31
5NHZERMnVZ3mcVYOrHt6tnrEsdXxntAEZn1qABk7z+wx9u9CCVabx1TJpD5+7LoKYaYxyjpj5njv
2oY9gymWe5vjoCmKzLN+YXF0P7YGIoQCqUvSGFfEOEEd/UavT5PsGxwtE9l1pWLKfrktlCoUnew9
2teX08SAchP0DFd4MG4o9gsBgUB7qL5vm5rncP33R1TOwUdd+nrpO4quyav/LukTed0SXus8E8Vz
lzM9Pv9+cjFVN7/t4a8i7prWk04MpWrG1Nr5RkIfHS17+zm5NQ4961Wv0IPR9E4zJUwDs7Hf59fo
hIzcTdpY65vh9ne8xgfOqn5JRbwnvy9AXC2K/i4a/uzOyuXBJ9TgxmQu766/kBRjdkzYi/HAp5nm
m1wDNylHspMB1FhI2qgqSOSWs+FMssLudpiNY0jGXFLSki12LGR937OOovfQ9JsB3KH6WD+su0+4
d8NNLC1s3SzvbI/GNW1ZI4WAsJ2NIqpEzX/sq+bL53VMCJKYX/JTkfNgQ+uMRBTeEFHLiWXpoWAu
1CvOpQOILtap/USVbxaPf4h2G5lq7Iczmg35xv5OM5AW8k+XRmg49drlU5c5oKOmMdtnC6jcHdnw
1gc/CqepPLzLi5q3AwpRc/yx6OJIEp/vWaS6bR1e4FIhcsR9aKdh4ZOxsgdsN0GIcmaOWbQZG7r3
Rj2OQqNQVImQD8OErURPzIHW+8Ck3K9JEfC2Gs4o/q13kyYp2cJvnaZZq9rJOKF69UxU4Kt6LOe3
gejTi7ritZpnm6k+9lIgYowbEpgIkPqPPPCdD5A9Zxf2H5xZw+9NDMfp0mUzNZGeLpKuBdPqOaRX
D9tOcVfJ4hqEKYguVbmHSY+i7+q0iuUwWIYYhKTdF3HJSJdSxYtjGytRrPwlOAMNq70M4dhRzp2U
GVPH3xjxB7petILsVsbqhHQCCchvt4tK15q/YhxWqaOQJhhy+Fy1u0EZ6PC2ZY/z1p3b2W6j8HhY
fzJRD0wVP038E0yHBvNlnnFXFwPZSEbvldm06pfKYQCnFs0MyHU6Bh8us/YfZnw/GUaM4XETe8lm
H5GQR3GbZvyoAoNcz1jG/IESGnN1EKr/DYIpk/jt1KznW1Iz1dmWhdc10+t7I5e3zZLxt7MEAxMN
XX/29f6Uc8v+6Pt35Ik9UxOxM0zeh2a2QqNykheAUJYw7LR1OjpO9RKaP66QEJcRuuKk/jFJCF3s
IbzQ1Qydth8o0Sxd2z7SnROSYRp0+2Bc/kDucuQ0jmFzU3noH6aQ4zwL7E4B4T7tOh5gCTVeQv5N
cuHYU3qExv75EQL2gTyOS0SemUXbY0FT2cxlDKnRm8r7mn/n9EWMfzkpt7Qy5y35/uiGOUDf75/T
KQL5wM8S9JWvEslkmygxbxthZLwt24RPvpCTybLkI4E/Gp9vcfQba+WYtP7MpJdgOTt3mkK4HbbQ
iGJA5Td287B8PCT3fTlRGne4ZKAlBeIxw36rL2+S1JlHMqFcjkMOVLcTAIq7sA/GbXSKUvWEzRxq
vyHRIDKiUjVmD9pu5FeYcPRapTquldPQRTt43uuMn+ogtxyEXOG7kP9PNkvKuaFyeIO7D/oCzxm+
lplAIZbzUDJcDrEvQ0v1trPk7VkOTopJLn1gLH3/moK3/KhxL8TLlUb9l8VoBNGG60oTj/v7l1n+
9499M35TKCSc90q9cOtGxN/6dZECD/KMKnw2BgyT6pdnM4SYdx+wTi+CGdTme4VPE9KAzQh9XE+u
jwR7HTbb8sXED+9QENwgkX0VpuPsQtP3v4eClfX0cg3yi4mUJmTZtWF8YogkjzsAFrFhPTG32HY1
zNyHTbaxj4oBi94hqRacR5eKEzUxGuuJ0zvcdq6mMocbcTd8F9qKq0aKenyQHncGEr56ntcEH7Ur
92XzX5G+SdulQ/XqQS+z2NX7JX4oSrET4fhrP0xvHFLSbr/IhHxRaklwpwr/vTNJ9bWTQApY06ws
z2UMbDBwbz6xJxlXzaKIzI9o8JfNt5wjoe7wJHRCurthVjFiyx6LCoNs1BG0C5/axpfJ4lGlEYpR
v+tyPsjaHCRIeKAOmTNG3OsojB5RjNkRMqOBeN7Rh49JMb8NkiibQeyY7FQXfxhnos6lVHlv4ITb
gQP83UXh+dzEmOjrkj2425uesKqKB6Wn2MvB59hrnrqZXtGJIOi/Y+52355KwPRCz5SifG6iyPmW
ahUzUU0oixjGcel1fdeOfKDGvEjkhnPdgJejTvCF0YQOp9PbtvSIyTZHDWDy7wDJFF8t434yzCBo
fI9REew6VK/SLfULLBvd2GaAS6+Z2aeAhRAaQhBYNB9bgsKx6UCKPX/S+VQ19hCrp+gV0yrRRqYY
n1lzQfP9GBDBhRBd14L6cG0LqVF7sNrsVDEztX83A1h/WBpFIJWzkerOg1kf51xHpTEwA5l8knzW
F1eZ7EKpYYU+VxwupqdolX8AyQFDzRO0MKmRw5Irg13zv2YsONI9JSQPZozRIDOrGDL9Nw6JWo8g
j3Iu/bWyvJlhadz/UOpct5/jvzE/1Qzt3Q+a1plIzV9hniPlEcBmOu0zOuM8xX9CBfYvWnzeXghs
WK7EV1cODkQRvrzKdoym+vLzw6lIxOyx0PhoXk9oVtFigLlssGAdMw7SRAw1jSWMAnot8nFA4p79
yeAoDbUJXNEnsvnuGR89HvQcZrfGKZJUDeGXVC14uu+7zq4ecldiN19PEBGJESm+pYQwbqRGYqCP
5CoDR7mOf8RFdqVM71fX9CJjU9v88rYzVgraS1cPGzzQurhNq2qHsjYQSu6/OPu0mzNxuOKn9xEX
sl2P1X5Y+RaVO0Hc+wtHIO0hs3upfqT0ZYx+jI0Ze9LaA4YABswvjHsDP55FatNL43fwG5g2Loe0
i+ubotboUiGbaye1D4irr7mrnqPJ7pPBfBHbTcpVHo9tz4bYgbXvU0Cpqv3c1ryzVPlduecYMHuo
bnpXnyzFRZlUGa73ZMJLbKnGabFFCknxTydEXaQP4j+e+7CUaqUjsK1o1JPm3QwKsiIfenAVu0/6
GEzmjXq9r8sxKs2BAsjCk1oVWLNecme+8p4uJU/xiOrIyciDb2lMQgS7MMloDycY2JQpOGWT7Z74
xKy4PZIwF/XZTo6H3+W2NDmp9XQ3jvWjWKWwfAnDzOhuBXQyvN8AoY5DQQkA/vt3gjQeEhHzOYpC
1RFtww/Gnq8lV6RssEYzKc2ng8/EDvOgSlQohGp+3+U4SEtBGPoMNVGRxaufmD5Z+00eWjCWqEa3
4wevTCllH3Md0z9OgV8Z0RlS6NZlrPCo8ZdewUB8M/TesSymvBFaLAsKfZbzfGoU2PawbY3AJe4L
f/7nTxc2tTYmF2VarfX1dsaoJBXTxTKRYZPR4La9/tL7qMFPOgoZO+modDtGaLddqzdrCZX0RCJM
O9N70fWmv+bzN7TZA9tfkQY5r0K0F1v/X6MXD1EQlrUVy+cvOzay9P9T6CwRSUSOO7exVQKQcJaV
n2ZynD/3t65L4644piY71wR4HQa5nFOSk1hvBg2HdTxUy/Ze/PuV7k1GiooEcUdtPV03TQ9BPhmS
LpCwwYnwtpKYzGI87jprfJJ58mW50fscN9875/hyqlinZ5mEe/O7290RrPbp3Ces8FpvGi4026GB
PuM+TD9oqJ6tjYnlJzSP5NqYQD7YNuDUaiTG1vdGdWDaZE9+jUch0LQ46VPMJF46g8fM5Gb4QQ9j
zrjEl0C/P3n60ooAKDPykibFqHdfjGVOVtYCqjZQxA3mCvCLA6RJcVg8W8E3RPRLOob/U/vy2T/1
43R4BvWnyR9aB4ZBo9SwUTB7ls+zkh0I/xYsnEhA1LyLjEuLc2iIKSiJRTktEbHRgUQ1SDey8C8X
9Op3p0gfd4eRymxFRKJR9H0iM7PpSB7dxRqRtpCdbqzCNLiCifZEKKeocH+AKy8Of5kSYWtTFMCh
FLZm6hxTIlxBX6lrbgTDJKqBUUe2O0wAKl/bj2hCloX6hw09TQILpgloQ5iJQElAmVVC1rKO24Wa
n/CyoSYgrKpSAFqLlNF0w5R7getRmVxf3KPgqcV+7IovjwwtrC3B2Gis3Q4AVE9izziGRVl/1OxI
IKJiP45lv53BmtNTIvWX1CWN5Td16gi3QiLGuqPjA9RrFo4/MFviXU1Wa1CI5L0kZZQkN+8ismUT
7ifLK9PEkFYaaCME9ngewVLYgcTRLMlrZVF/WRUy7LubW2W9EESQfwmeZ1t7SBNC0IQb45JfC08C
iuNxmIr1nyszmG/hDGlOgQK4t876QB0xyPONw0Bwu+D+balvZAUQRRuOqimLv+e8YHFp6jXgVGOL
A/iOGtIYjuMcTDbH+AIAR6p05jeORrd6SazaXqGFF46l2xNKRXe/MsGWyylyjY+ebrQmU3BLbov/
tdjOIcw7UfYPhdUx01CctIB+rMWx1CP5cicL2TAuDA8gwAGdb0NkDV093lV6Id0ciIsJbtb2qjpu
PJBzGE/AJP/bTwajHyKNgA4pYcZeFTIzDazJyU0zyzQCEtVdWViLneDlIvkXLd2ELEIOQEOKPeDW
lMAsTh7lmxVoTMj1J/+IylY1uV6ftzXioA/oHvX/TG/sfKPDCvP1FztKZYlz/5TyvXcHLv21I8He
JUrD5bJtjwCplL2inQIjDi/9T+nL26qyzQDm5vp0h/EBfs6/dQNPESWP//kFFT6F0f+qUnZvBE5/
mu1t1xhJbBn67dLgaekO4gaXQG8jroaapt+TdRRsnDYhU/A8caqYFO1wOw1shZS+JxZRfMQs5ZWX
Otls/c+Hi+aRM1qlqqujjMIg7ESy4M3wScXrYjvuOO7UQ/XUUTmwZg33/4K2kTFpLI2lcMZG9VNI
PZMkDmHLjfxGybXPW1+QIv6eDZ2mmpGgXlMM7yTzfz4iuBZoW6rcjwnDG3wuKVTiuU2zrEZxnhwl
Q0ChsEQdGYE5efxuveD30yu/CIJV7bNBFGIyFvEBYkcjXBzFDAhBaLWna2LYrDfOqdMcoYNx4xGe
vGXgnbOW3SBJDMnDJSmLNXonzFGyhOJ94YTaXiBOAY4O8fMIn/05oVFCYpOt+Qm5aswOWxCg/ay5
BWw3BAiyttC1D8A5CejS8KO8PNt2iVSzM2VQvDd2C7sgU0ljchKW8UFByShKZSWYEQIqyWENauYl
b9fjS8WN+Bn1CjP6mUDtMh2H9ZyHsTyGhJB3M4+toF6gGUdl+N0HX044Do6eC32lwmdLqmFFJ3+v
j0sZngHSltHH+4Hs3MQScR7vj8Gq7bIQc7hBz8CqOCHCTyKuH0YzgZiP6gyyW7+BIaKi2AFr0hrs
2iJXkr31yLVybjjQ7rc0gN4OSK2HnRPTh74k1qNiilFlX8bADhl6CWy+803pgdUWp3+GCiNOgYLH
NC4XcP+iLrkVCqPZWvzwwTWos+L4x/tGxl3PotZF3LD9ECDqxdjZKuPex4yowyV6VBSXBycXc4Qo
O8ca3c+XtE8KgxVT1QF/FXI=
`pragma protect end_protected


endmodule
