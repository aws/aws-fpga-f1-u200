// Amazon FPGA Hardware Development Kit
//
// Copyright Amazon.com, Inc. or its affiliates. All Rights Reserved.
// SPDX-License-Identifier: Apache-2.0

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Xj78u+crC0DVwcb6TXHWKv4w0HzS32NHDZyGOH8cqWQOwvNROgoHijIoIBayPYeih9IOmLmoI4It
LVnXCSxJ2/DeOebRH1OEKZPeHqNW9rI6qdksXtBr+yibD1ivz6p4tDLUi9RQCSl1szINoo3EECxV
i9UBB174TeK1yKcv45fFdqDMXJJi+8aj6V5pQEQvV+UIZxIeqygK+lAul2b0nscPEqV+H3xfjEW9
u+9IIhD7n51Hw6bwWqYYKjJze4vqm0voTAfPB1GkczbxuzElLZecvIu/uRBq4eJrMv/VIPiQ1mfK
J60fdHXRBXaofmt+drl1gB3bV99DQPzBpt3xrw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
na2HRJ8to9+QolGwJXsQPBynVTAM6r0OFOXwAknXLKC/+essXWwY7Pn2Fnj0/cUC9HddU5PRr+Nn
KCpVJYCMLnmWH60kztZsSj2RYgCq39FpKfwUzTSRztH3CT7g6rBmzSVQMr7JpSZ3ZugN/uHjY1u/
irEUyx7b98ZXrwTn8kM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
IWNkpf/IPFwtENrGYBNqA/+hgSM9cVrSRlzNRD/WDjKwqHQ5adCkXIAY6LIdXDXNT72c6Pe19W5x
QvEQRnviKVQShk4XMXHT/WMuUJe46A66FABcO5BDGBn1TFH+KP9denQXGjN6kYYCiQ/tXSyWXehj
b0d3ucAWNDJtkiEGaG8=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
JnK9rXuV3P5G9YUNo3fU8uKlaqn/8z7mHKg8UXtvOxeQYxCVTd7U9Z3e0jvI7tGp0FBigYHEdLDl
EWo+C5vS/Q==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2256)
`pragma protect data_block
VxVHqqYFpHvKKNAdD+yGkDdKDS0OSsZVxs3kpUU2WRtpJYEIEE63mRk1mMErB6Zdq1tUKd2xtsDc
ET8+bUtzFgSmdwSq1BbTA9HtgmAxdbFZhwnPUq1kGxs1oVfu4pohBJfVuawS5DcuzSKVAq7KKR1L
vXV145mx5NU2hXgrpIxGjCAJqV/orV51YYzydWIPMj5qHzJVDz3MmgZomftepbTjeq0CjCVjF0Dm
XGmAaq3iVww5GMjxVVYNXA+wLv29zREfktpYrlBsX6oVRR4btzDYC/4gaxWhmvf/jY1sgz+rWqt+
GyPWRumacsZgnwyqb3/IwdXFaDGj/Z8Ii5hEAMa30DQJBQtEUQWsBY6xXw8OkrHtw+HCM+5wx3Tg
Y0FNM2AKmUESzyrLtlkJIXlefc/vLloPvbWgqltH9wRHIx7QEamE+vG+KxynRmnCPwPv0Btm3Srk
++AOFQGKUgHarYaQfjCjTzEn+I/YxKClM4bb5y8h9Wgpb7T6dHgAjEbcjHVD9fYPWuIf2hRCIhAG
a7/LlI4npTsvBITbum7f/+ZYGDuiUkc7LN5qDyut5x02MP/a1OCA0z9hrb+aDAq4MTY8BP/ek0ZR
sJlNtvDMKpmAvCaVtGnL2pO/VozEw6JqU2Ialm/NosuCjjrzNPSbwmR4bvnHY271E0jHFWYzJEaF
tOlu6a58hLU8SbzGi6sXK7P0JIIYCQmlOPJnZTMu1TfECofXLvEdymp8muXyfp0g0yybjfvqtNBX
Nu4GN7M4tovir5beq4LED7BKe6nllbft74zbZqDLtZTT+FxsGHIkw/Et9AgPxQtQo2GUZeGieGvV
J+4C/wsdoFgW74Nvd241yQXbvWAJBDOxozNPrO5YpQAOvqpPknt69hrqK1n83o6TwL0UA8rcYNBa
XtxvOboiGoeQCHcvCU1KfTxZPjDjY6wb8XS3l/wRvCRjyzj5gCOFF83QW92lYM9aqRL7k8enZSRv
ZqoQy4+GF/hIjEoY6Il2kXg4JOSdRL7RSGEq+ZKtL+7ovSoqb3n95HL21T1vO/xegiwqKSCxgs4y
ilrIVc0CdkofKc0V4n2hB4ch+sU5DefslCBQYokvUob/RGl0JqETKWvbG5NlFxTRHx6Fz0rJQawQ
YwKARD7JHtqODY07n1GZZBqCeBQhEkgLN8kMJPN9KJ6Jgp6DdgR+fF1o3kAsi9dR0ZL3sPoVnvHC
bwSWMzFoYQsPin2PBXcIvdDIT1iin35PrNv5muz2uICh5RkAWNMoj/xuZkdPyVHzYwOXQrkBvOkM
vU5r2riX3N6yUfo2U3nFLjzkrq0MJ28Zf4p+Ya8YMGlSazxpTNMyznZkivE1FicgumwtDMYjvzUY
MA4PK4F+IGHI3+cXap0jr3RfImWw4OJGeqtrosMIv6Sab/9S04lCMYH6jK4OsDKnS5HSm/fme1Uf
D6WVVQK4hfx7oQhv0Eyg4Qm0rrdapkqEsce8uNJeCX8H/ROlKakLATEieUJRRR7ViwRFm/GrKcI+
zs71oOM7dTwOjQ1ryW8Z8zE5fW3w4BfHTGLWt6jGBALHELFHnI4etGWNwCP2QjuQCRdO5boHV0AC
PZyh/tfmdaKK2Ir+kwT1MN8PlBka5dZeeJj193Kar6+A9ZD0Lvz58y/wMrN4mKjN3OJVr/lc/zMy
/vEUIdFXqQ/tcGxLWv0laJhNLC1bCGXYqISbKBI8ClXhHt9e75xih0MLbuvGx/pcKW4TCMXEP3Yo
JD3RaE/qtGgfZQw4gnxKlaHGz/h1rUEHpNrYlUm3Vu/zTxH3VExjkN0ViHXrD9HqMDdOJ3bfv61+
OZ1qlx+qIWkhkNwyxY+BlHu9RdOJ9RAECWjbqr1TUHUAbz2DKjv72R4SfZrwFJMv1o3KnBALkOMJ
jZ6Dfq+zu9mBo34cBdCrHEzNVOEa5WHxg6Gukud64lmXb0lFFRKrkFfvZ1XPUfbOLHPRbPECjVwJ
aXjbzFxDBEiOCZ5UwFdwdDs0yHjgE4xyUhVmYXiMVgfwUcPBeRWsSGb1AYNEswvHGWbFWjyzqxID
JYR8pYM+wVv0E5rzpbtRwWGwN0IFEr1l+7O4XYbiEseXs/Lf+RTmFmKWSlWAFOjr+QvUeHa/PZ8S
BeKNQdbtDisPNnVwc+vfZFpJXtfxVz/gSqajXwE+HY/p+mMiD5fjFAjahm4OPjFvSrJhkQJoL5Yd
raJ++c6C9AKKikA55u2WHREW6WH9mWCVuBIhNHq7QRpUH8TIBbra4V5TAQWTnD6uhFQINm5qeWl4
tGaOx+AKUJ70O7gVtWZPq/r78yz6b8VWZ105StGuRzCZU0kkcsMr15XuPv2HpxjAv+Xi/TaNsoW3
xZYbBeDYq7u/alO8lzqLDCHCwSHtZUgGIeEbChxNPeIiOPuqoWT3VBfxrouTNfSdhBEDKYUoXNnT
B0Zs6JANeoK/zLQ3tVzC9zgvNXnh/OSrr+vs0XRSber00mcZ1iUNhWCl9xhEow8gocT58OyQwHfE
fkSBX/0CluqxWGNxh1aqpKKEjlEL8/jb5Sv1JQJW3HKtnpsiiP/i4VM61VJgirWPaO6k2oYIiDyI
vrq+UYZVpb3zgE+BMyLhMz7zPIVdBguSm3exTEkzOhA0GOZHaJfE8NqiCe5l0d/p2H4HL2QyuHuQ
5XiS48QEF5aEFwvc9KnlrPCC7RZS0HwNT06sCA9uJ59sONtVD3kyed4897dbE1lXlR9mZyrENHmE
5dzPs0vQQeSd7T9brC2V1t5rQWFplSJtPetvJZlLXaJmknN7JCZ43QLN4XvZ+UhodJflPIfjeEmt
ICg9I4Csa0NWp5JqcLt1gy/3SXuDlNz/DtNLT7Lc8hUmVUO83XLBhUM4w+OXVHjMx2wRAqKvE40G
+ddP937J/wZY+x/ergL4Z+UH2DYwFQl2kdeWFJYVdUjvQoUeDQRhe1RUUnVDed0sXLlowLuzpMHx
/24A9scg5xGXq7uKw051Pd5OawGd04m1GRAgGRpex3A5
`pragma protect end_protected
